library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity texture_rom is
port(

	--clk : in std_logic;
	tex_addr : in unsigned (13 downto 0);
--	side_in  : in std_logic;
--	texNum_in : in unsigned (3 downto 0);
--	texNum2_in : in unsigned (3 downto 0);
--	bool_in   : in std_logic;
--	
--	side_out  : out std_logic;
--	texNum_out : out unsigned (3 downto 0);
--	texNum2_out : out unsigned (3 downto 0);
--	bool_out   : out std_logic;
	tex_data : out unsigned (23 downto 0)


);
end texture_rom;


architecture rtl of texture_rom is

type rom_type is array(0 to 16383) of unsigned(23 downto 0);
--constant ROM: rom_type := (
--
----Red Brick texture MSB = 00
--
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
--x"49",x"c0",x"a0",x"a0",x"a0",x"c0",x"80",x"a0",x"c0",x"80",x"a0",x"a0",x"60",x"25",x"49",x"49",x"c0",x"a0",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"25",
--x"49",x"c0",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"80",x"60",x"60",x"25",x"49",x"49",x"c0",x"a0",x"80",x"80",x"a0",x"80",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"a0",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"60",x"60",x"25",
--x"49",x"c0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"25",
--x"49",x"a0",x"a0",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"80",x"a0",x"80",x"80",x"80",x"a0",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"60",x"80",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"a0",x"80",x"40",x"25",
--x"49",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"80",x"60",x"40",x"40",x"25",x"49",x"49",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"80",x"60",x"60",x"a0",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"25",
--x"49",x"a0",x"a0",x"60",x"80",x"40",x"60",x"60",x"40",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"80",x"80",x"60",x"60",x"40",x"80",x"60",x"60",x"80",x"60",x"40",x"60",x"80",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"40",x"60",x"60",x"40",x"80",x"40",x"60",x"40",x"80",x"40",x"60",x"40",x"80",x"60",x"40",x"60",x"80",x"60",x"80",x"40",x"25",
--x"49",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",
--x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
--x"a0",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"40",x"49",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"80",x"80",x"a0",x"80",x"a0",x"80",x"60",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",
--x"80",x"a0",x"80",x"a0",x"60",x"80",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"80",x"60",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"49",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",
--x"60",x"a0",x"a0",x"80",x"80",x"60",x"a0",x"60",x"80",x"80",x"80",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"a0",x"80",x"60",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"a0",x"60",
--x"a0",x"80",x"80",x"a0",x"80",x"60",x"60",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"60",x"a0",x"60",x"80",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"80",x"40",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",
--x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"80",x"40",x"80",x"60",x"60",x"a0",x"80",x"60",x"40",x"60",x"a0",x"60",x"80",x"40",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"24",x"49",x"49",x"a0",x"60",x"a0",x"a0",x"40",x"a0",x"60",x"80",
--x"60",x"a0",x"60",x"60",x"40",x"60",x"60",x"80",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"80",x"60",x"80",x"80",x"40",x"80",x"60",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"40",x"24",x"49",x"49",x"a0",x"a0",x"60",x"60",x"40",x"60",x"80",x"60",
--x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"49",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"24",x"49",x"49",x"a0",x"60",x"40",x"60",x"40",x"40",x"60",x"40",
--x"25",x"25",x"25",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
--x"49",x"c0",x"80",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"c0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"a0",x"80",x"80",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"40",x"25",
--x"49",x"c0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"60",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"25",x"49",x"6d",x"c0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"40",x"25",
--x"49",x"a0",x"60",x"a0",x"a0",x"60",x"80",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"a0",x"80",x"60",x"60",x"a0",x"60",x"40",x"25",x"49",x"6d",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"60",x"40",x"25",
--x"49",x"a0",x"a0",x"80",x"a0",x"40",x"a0",x"40",x"60",x"80",x"a0",x"80",x"60",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"40",x"40",x"25",x"49",x"6d",x"c0",x"60",x"a0",x"60",x"80",x"80",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"60",x"40",x"25",
--x"49",x"a0",x"60",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"40",x"60",x"60",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"a0",x"80",x"60",x"40",x"60",x"80",x"60",x"40",x"25",
--x"49",x"a0",x"a0",x"60",x"60",x"60",x"60",x"40",x"60",x"40",x"60",x"60",x"80",x"60",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"80",x"60",x"80",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"40",x"a0",x"40",x"60",x"a0",x"40",x"60",x"80",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"60",x"60",x"40",x"25",
--x"49",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"25",
--x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",
--x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",
--x"a0",x"60",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"80",x"60",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"a0",x"60",x"80",x"80",x"80",x"60",x"80",x"60",x"80",x"80",x"60",
--x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"40",x"a0",x"40",x"80",x"80",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"49",x"49",x"6d",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",
--x"a0",x"80",x"60",x"a0",x"80",x"a0",x"80",x"60",x"80",x"60",x"40",x"49",x"49",x"49",x"c0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"80",x"80",x"60",x"80",x"a0",x"60",x"40",x"49",x"49",x"6d",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",
--x"a0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"49",x"49",x"49",x"c0",x"60",x"a0",x"60",x"40",x"80",x"a0",x"60",x"80",x"80",x"a0",x"80",x"a0",x"60",x"80",x"40",x"60",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"80",x"60",x"a0",x"60",x"a0",x"60",x"80",x"80",x"a0",x"60",x"80",x"a0",x"60",
--x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"40",x"49",x"49",x"49",x"80",x"60",x"a0",x"a0",x"40",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"80",x"60",x"a0",x"80",x"60",x"80",x"60",x"80",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"40",x"a0",x"60",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"a0",x"60",
--x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",
--x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
--x"49",x"c0",x"a0",x"80",x"80",x"a0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"40",x"a0",x"80",x"40",x"80",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"a0",x"40",x"25",
--x"49",x"c0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"80",x"60",x"a0",x"60",x"80",x"40",x"a0",x"80",x"60",x"a0",x"40",x"80",x"80",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"60",x"80",x"60",x"60",x"40",x"80",x"40",x"80",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"40",x"25",
--x"49",x"c0",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"80",x"80",x"40",x"60",x"a0",x"40",x"80",x"40",x"80",x"60",x"80",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"60",x"60",x"80",x"a0",x"60",x"40",x"a0",x"60",x"40",x"80",x"a0",x"40",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"40",x"25",
--x"49",x"c0",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"80",x"a0",x"60",x"a0",x"40",x"80",x"a0",x"40",x"80",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"60",x"40",x"80",x"60",x"a0",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"a0",x"80",x"a0",x"40",x"25",
--x"49",x"c0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"80",x"60",x"a0",x"40",x"24",x"49",x"49",x"c0",x"a0",x"60",x"60",x"a0",x"60",x"60",x"40",x"a0",x"40",x"a0",x"40",x"80",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"60",x"a0",x"60",x"80",x"80",x"60",x"60",x"40",x"25",
--x"49",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"80",x"60",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"60",x"40",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"40",x"24",x"49",x"49",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"40",x"60",x"a0",x"60",x"40",x"80",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"40",x"25",
--x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",
--x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"49",x"25",x"25",x"24",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",
--x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",
--x"60",x"a0",x"40",x"a0",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"a0",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"60",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",
--x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"40",x"60",x"60",x"80",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"a0",x"60",x"60",x"40",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"80",x"40",x"a0",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"40",
--x"a0",x"60",x"40",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"40",x"a0",x"80",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"60",x"60",x"a0",x"60",x"60",x"60",x"a0",x"40",x"a0",x"40",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"40",x"80",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"60",x"a0",x"a0",x"80",x"60",x"80",x"60",x"60",x"60",x"80",
--x"60",x"80",x"40",x"80",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"60",x"60",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"40",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"40",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"40",x"a0",x"80",x"60",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",
--x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"80",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"40",x"a0",x"a0",x"60",x"a0",x"60",x"60",x"80",x"40",x"60",x"40",x"a0",x"60",x"a0",x"60",x"60",x"60",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"60",x"40",x"a0",x"60",x"a0",
--x"60",x"a0",x"60",x"60",x"60",x"80",x"80",x"60",x"80",x"60",x"60",x"40",x"a0",x"60",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"40",x"a0",x"60",x"a0",x"60",x"60",x"60",x"80",x"40",x"80",x"60",x"80",x"40",x"a0",x"60",x"60",x"a0",x"80",x"60",x"a0",x"40",x"a0",x"40",x"80",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"40",x"60",x"40",x"a0",x"60",x"a0",x"60",x"40",x"60",x"a0",x"40",
--x"60",x"80",x"40",x"a0",x"60",x"60",x"80",x"60",x"60",x"60",x"a0",x"40",x"a0",x"60",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"40",x"60",x"a0",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",x"60",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"80",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"40",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",
--x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"24",x"49",x"49",x"a0",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
--x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--
----Blue Stone Texture MSB = 01
--
--x"49",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"49",x"49",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"25",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",
--x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
--x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",
--x"00",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
--x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",
--x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"24",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
--x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",
--x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
--x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
--x"00",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
--x"00",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"00",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"00",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"00",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"03",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
--x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",
--x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",
--x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
--x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
--x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
--x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
--x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",
--x"24",x"24",x"24",x"24",x"24",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"00",x"24",x"02",x"01",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"00",x"24",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"03",x"4b",x"03",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"01",x"01",x"02",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
--x"49",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--
----Wood Texture MSB = 10
--
--x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
--x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",
--x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",
--x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
--x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
--
----Mossy Texture MSB = 11
--
--x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"d4",x"d4",x"d4",x"d4",x"d4",x"db",x"db",x"db",x"db",x"db",x"db",x"b4",x"b4",x"b4",x"db",x"24",x"49",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"d4",x"d4",x"d4",x"6d",x"92",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"da",x"b4",x"b4",x"b4",x"b4",x"92",x"b6",x"d4",x"d4",x"da",x"b6",x"b6",x"d4",x"d4",x"92",x"24",x"49",x"92",x"b6",x"b6",x"92",x"d4",x"6d",x"d4",x"90",x"90",x"90",x"6c",x"49",x"49",x"49",x"24",x"49",x"6d",x"90",x"90",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"24",x"49",x"49",x"db",x"da",x"b4",x"b4",x"b4",x"6c",x"92",x"d4",x"d4",x"90",x"b6",x"b6",x"b6",x"90",x"b4",x"6d",x"24",x"49",x"b6",x"db",x"b6",x"92",x"6d",x"d4",x"6d",x"6c",x"90",x"6c",x"49",x"6d",x"49",x"49",x"24",x"49",x"90",x"d4",x"d8",x"90",x"6c",x"92",x"b6",x"b6",x"d4",x"d4",x"d4",x"6d",x"6d",x"d4",x"d4",x"92",x"92",x"92",x"92",
--x"da",x"b6",x"b4",x"b6",x"b6",x"b6",x"92",x"92",x"24",x"49",x"49",x"db",x"da",x"90",x"90",x"90",x"6c",x"92",x"d4",x"90",x"b6",x"b6",x"92",x"92",x"92",x"90",x"49",x"24",x"49",x"92",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"6d",x"90",x"6c",x"49",x"6d",x"49",x"49",x"24",x"49",x"90",x"d8",x"b4",x"6c",x"6d",x"6d",x"b6",x"db",x"d4",x"d8",x"d8",x"49",x"6d",x"d4",x"d4",x"90",x"6d",x"da",x"da",
--x"b6",x"b6",x"b4",x"b4",x"49",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"db",x"b6",x"90",x"90",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"90",x"92",x"6d",x"92",x"90",x"49",x"24",x"49",x"49",x"b6",x"d4",x"90",x"b6",x"92",x"92",x"6d",x"48",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"90",x"d8",x"6c",x"6d",x"92",x"b6",x"d8",x"d4",x"6d",x"90",x"90",x"49",x"6d",x"90",x"90",x"6c",x"49",x"92",x"92",
--x"b6",x"92",x"6c",x"49",x"92",x"92",x"92",x"6d",x"24",x"49",x"49",x"db",x"da",x"90",x"6c",x"6c",x"6d",x"b6",x"92",x"92",x"92",x"90",x"92",x"92",x"6d",x"92",x"49",x"24",x"49",x"49",x"6d",x"90",x"90",x"b4",x"92",x"b6",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"90",x"90",x"6c",x"6d",x"6d",x"d4",x"d4",x"d4",x"6d",x"6c",x"90",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"b4",x"6d",
--x"b6",x"b6",x"6d",x"92",x"b6",x"92",x"6d",x"49",x"24",x"49",x"49",x"db",x"da",x"92",x"6d",x"6d",x"92",x"b6",x"92",x"da",x"6d",x"90",x"92",x"b6",x"92",x"92",x"49",x"24",x"49",x"49",x"6d",x"92",x"b6",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"49",x"49",x"49",x"25",x"49",x"90",x"6c",x"6d",x"92",x"92",x"6d",x"d4",x"6d",x"6d",x"6c",x"6c",x"49",x"6d",x"6d",x"92",x"6d",x"6d",x"90",x"6d",
--x"92",x"b6",x"b6",x"6d",x"6d",x"92",x"49",x"49",x"24",x"25",x"49",x"db",x"b6",x"b6",x"92",x"6d",x"92",x"d4",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"92",x"49",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"6d",x"92",x"6d",x"b6",x"b6",x"6d",x"92",x"b6",x"6d",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"6d",x"6d",
--x"92",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"25",x"49",x"db",x"db",x"b6",x"6d",x"92",x"6d",x"d4",x"b4",x"6d",x"92",x"92",x"92",x"b6",x"92",x"92",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"90",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"92",
--x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"db",x"db",x"92",x"6d",x"92",x"92",x"d4",x"90",x"6d",x"b6",x"92",x"b6",x"92",x"b6",x"92",x"49",x"25",x"24",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"90",x"49",x"92",x"b6",x"d8",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"6d",
--x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"db",x"b6",x"92",x"6d",x"d4",x"b4",x"90",x"6d",x"92",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"6c",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"90",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"49",x"49",x"92",x"db",x"da",x"92",x"6d",x"92",x"90",x"6d",x"92",x"92",x"b6",x"6d",x"92",x"90",x"92",x"49",x"49",x"24",x"49",x"49",x"6d",x"b6",x"fc",x"fc",x"db",x"db",x"db",x"da",x"da",x"db",x"d4",x"6c",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",
--x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"6d",x"b6",x"da",x"92",x"b6",x"92",x"92",x"92",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"25",x"49",x"b6",x"fc",x"d4",x"90",x"92",x"92",x"b6",x"92",x"b6",x"90",x"6d",x"48",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"da",x"b6",x"92",x"b6",x"92",x"6d",x"92",x"92",x"6d",x"92",x"b6",x"90",x"49",x"49",x"49",x"24",x"25",x"49",x"b6",x"d4",x"90",x"6d",x"b6",x"92",x"d8",x"d8",x"92",x"90",x"49",x"6c",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"b6",x"92",x"d4",x"90",x"6d",x"b6",x"92",x"b6",x"92",x"6c",x"49",x"6d",x"49",x"24",x"25",x"49",x"b6",x"d8",x"90",x"6d",x"92",x"d4",x"d8",x"6d",x"92",x"90",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"25",x"24",x"49",x"49",x"b6",x"b6",x"90",x"92",x"90",x"90",x"b6",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"d8",x"d8",x"6d",x"6d",x"b6",x"d8",x"d8",x"6d",x"92",x"6c",x"49",x"49",x"49",x"49",x"d8",x"b4",x"b4",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
--x"da",x"d4",x"b4",x"db",x"db",x"d4",x"90",x"6d",x"6d",x"49",x"24",x"49",x"49",x"92",x"b6",x"6c",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"24",x"24",x"49",x"d8",x"6d",x"92",x"6d",x"92",x"90",x"6c",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"b4",x"b4",x"90",x"6d",x"25",x"49",x"6d",x"b6",x"d4",x"d4",x"d4",x"db",x"b4",x"b6",x"b6",x"d4",x"d4",x"d4",x"db",
--x"d4",x"b4",x"90",x"b4",x"b4",x"90",x"6c",x"49",x"6d",x"49",x"24",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"92",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"49",x"6d",x"92",x"6d",x"92",x"d8",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"90",x"90",x"49",x"6d",x"24",x"49",x"92",x"d4",x"d4",x"d4",x"6d",x"d8",x"90",x"6d",x"b6",x"d4",x"90",x"90",x"6d",
--x"b4",x"90",x"b6",x"b4",x"90",x"90",x"6c",x"49",x"6d",x"49",x"24",x"49",x"49",x"49",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"25",x"24",x"24",x"25",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"90",x"90",x"6d",x"49",x"24",x"49",x"92",x"d4",x"d4",x"6d",x"92",x"90",x"90",x"6d",x"92",x"d4",x"90",x"90",x"6d",
--x"90",x"b6",x"92",x"b4",x"90",x"6c",x"6c",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"90",x"92",x"49",x"24",x"49",x"92",x"b6",x"6d",x"92",x"92",x"90",x"6d",x"6d",x"b6",x"d4",x"90",x"90",x"92",
--x"b6",x"92",x"b6",x"b4",x"6c",x"49",x"49",x"92",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"92",x"b6",x"92",x"b6",x"49",x"24",x"49",x"92",x"b6",x"92",x"b6",x"92",x"b6",x"6d",x"b6",x"6d",x"b6",x"90",x"6c",x"6d",
--x"92",x"b6",x"6d",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"6d",x"49",x"25",x"49",x"6d",x"b6",x"db",x"b6",x"b6",x"6d",x"24",x"49",x"92",x"92",x"b6",x"d8",x"92",x"92",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"92",
--x"92",x"d4",x"90",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"92",x"d4",x"d4",x"b4",x"90",x"92",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"90",x"d4",x"d4",x"d4",x"b4",x"da",x"db",x"db",x"db",x"d4",x"d4",x"d4",x"d4",x"b4",x"90",x"90",x"24",x"49",x"6d",x"db",x"b6",x"db",x"b6",x"6d",x"24",x"49",x"6d",x"92",x"b6",x"92",x"92",x"b6",x"92",x"d8",x"92",x"6d",x"b6",x"92",x"b6",
--x"92",x"90",x"90",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"d4",x"b4",x"b4",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"90",x"d4",x"b4",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"90",x"6d",x"90",x"90",x"90",x"90",x"6c",x"24",x"49",x"92",x"db",x"b6",x"b6",x"b6",x"d8",x"24",x"49",x"d8",x"b6",x"92",x"b6",x"92",x"d8",x"d8",x"6d",x"b6",x"92",x"92",x"b6",x"92",
--x"92",x"90",x"92",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"49",x"b4",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"92",x"db",x"92",x"92",x"90",x"92",x"d4",x"b6",x"92",x"92",x"6d",x"b6",x"90",x"6d",x"90",x"6c",x"48",x"24",x"49",x"92",x"d8",x"92",x"92",x"b6",x"90",x"24",x"49",x"90",x"48",x"6d",x"6d",x"d8",x"b4",x"90",x"6c",x"48",x"6d",x"6d",x"49",x"6d",
--x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b4",x"90",x"6d",x"6d",x"92",x"90",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"d8",x"b6",x"92",x"d4",x"90",x"92",x"d4",x"d4",x"b6",x"92",x"90",x"b6",x"90",x"6d",x"48",x"24",x"49",x"92",x"b4",x"6d",x"92",x"b6",x"6c",x"24",x"49",x"48",x"49",x"49",x"49",x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"b4",x"90",x"6d",x"92",x"92",x"6d",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"d4",x"b6",x"d4",x"90",x"6d",x"92",x"d4",x"90",x"92",x"b6",x"92",x"92",x"6d",x"6d",x"48",x"24",x"49",x"92",x"6d",x"92",x"b6",x"db",x"48",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",
--x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"49",x"49",x"49",x"db",x"6d",x"92",x"b6",x"90",x"92",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"b4",x"92",x"d4",x"6c",x"6d",x"b6",x"92",x"b6",x"92",x"6d",x"b4",x"90",x"6d",x"6d",x"48",x"24",x"49",x"d8",x"db",x"b6",x"db",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",
--x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"24",x"db",x"92",x"92",x"b6",x"90",x"92",x"6d",x"6d",x"6d",x"48",x"24",x"49",x"92",x"db",x"b4",x"b6",x"90",x"6c",x"6d",x"92",x"6d",x"92",x"b6",x"92",x"b4",x"90",x"6d",x"49",x"48",x"24",x"49",x"b4",x"db",x"b6",x"b6",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"6d",x"92",x"b6",x"b4",x"b4",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"24",x"db",x"b6",x"da",x"92",x"6c",x"b6",x"92",x"6d",x"6d",x"48",x"24",x"49",x"92",x"db",x"b6",x"d4",x"90",x"6c",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"b4",x"90",x"92",x"49",x"48",x"24",x"6c",x"90",x"db",x"b6",x"b6",x"b4",x"49",x"24",x"49",x"6c",x"90",x"90",x"90",x"b4",x"b4",x"90",x"90",x"49",x"49",x"49",x"49",x"49",
--x"6d",x"b6",x"b4",x"b4",x"90",x"6d",x"b6",x"b6",x"b6",x"b6",x"49",x"24",x"db",x"b6",x"92",x"b6",x"6d",x"92",x"6d",x"92",x"6d",x"48",x"24",x"49",x"6d",x"92",x"d4",x"90",x"6c",x"6d",x"6d",x"b6",x"92",x"92",x"6d",x"92",x"b4",x"90",x"6d",x"49",x"48",x"24",x"49",x"90",x"db",x"db",x"b4",x"90",x"49",x"24",x"49",x"6d",x"90",x"6c",x"90",x"90",x"90",x"b4",x"b4",x"b4",x"90",x"92",x"49",x"49",
--x"6d",x"b4",x"90",x"90",x"6d",x"92",x"b6",x"b4",x"b4",x"6d",x"6d",x"24",x"db",x"da",x"b6",x"92",x"b6",x"90",x"92",x"b6",x"6d",x"48",x"24",x"49",x"49",x"92",x"90",x"6c",x"6d",x"6d",x"92",x"92",x"b6",x"6d",x"92",x"6d",x"b4",x"90",x"6d",x"49",x"49",x"24",x"49",x"90",x"db",x"b6",x"b4",x"6c",x"49",x"24",x"49",x"92",x"6d",x"6d",x"90",x"90",x"90",x"90",x"6c",x"6c",x"6c",x"6d",x"49",x"49",
--x"6d",x"b4",x"90",x"6d",x"6d",x"b6",x"6d",x"b4",x"90",x"6d",x"6d",x"24",x"db",x"92",x"92",x"92",x"b6",x"92",x"92",x"6d",x"6d",x"48",x"24",x"25",x"49",x"b6",x"db",x"b6",x"d4",x"d4",x"90",x"92",x"6d",x"6d",x"6d",x"6d",x"b4",x"90",x"6d",x"49",x"25",x"24",x"6c",x"92",x"da",x"b6",x"b4",x"48",x"49",x"24",x"49",x"db",x"b6",x"b6",x"90",x"6c",x"6d",x"6d",x"48",x"6d",x"6d",x"6d",x"49",x"49",
--x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"92",x"b4",x"6c",x"6d",x"49",x"24",x"db",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"48",x"24",x"25",x"49",x"92",x"db",x"b6",x"d4",x"90",x"6c",x"6d",x"92",x"92",x"92",x"b6",x"90",x"90",x"6d",x"49",x"24",x"24",x"90",x"92",x"da",x"b6",x"90",x"6c",x"48",x"24",x"49",x"da",x"b6",x"92",x"90",x"6c",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"49",x"49",
--x"6d",x"b6",x"b6",x"92",x"b6",x"b6",x"b4",x"90",x"6c",x"6d",x"49",x"24",x"db",x"b6",x"6d",x"92",x"d4",x"b4",x"6d",x"92",x"6d",x"48",x"24",x"24",x"49",x"6d",x"da",x"b6",x"90",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"b4",x"90",x"6d",x"6d",x"49",x"24",x"24",x"49",x"92",x"da",x"92",x"6c",x"48",x"48",x"24",x"49",x"b6",x"b6",x"b6",x"90",x"6c",x"6d",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",
--x"6d",x"db",x"92",x"b6",x"92",x"92",x"90",x"6c",x"6c",x"6d",x"49",x"24",x"b6",x"db",x"92",x"92",x"b4",x"90",x"92",x"b6",x"6d",x"48",x"48",x"24",x"49",x"49",x"b6",x"db",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"90",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"49",x"49",x"6d",x"b6",x"6d",x"6c",x"48",x"48",x"49",x"49",x"b6",x"b6",x"92",x"90",x"90",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"49",x"49",
--x"6d",x"db",x"b6",x"b6",x"92",x"92",x"6c",x"6c",x"6d",x"6d",x"49",x"24",x"b6",x"db",x"6d",x"b6",x"92",x"92",x"92",x"92",x"6d",x"48",x"48",x"24",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"6d",x"db",x"b6",x"92",x"b4",x"90",x"92",x"6d",x"92",x"92",x"49",x"24",x"92",x"db",x"b6",x"6d",x"b6",x"b6",x"6d",x"92",x"6d",x"49",x"48",x"24",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"48",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",
--x"6d",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b4",x"90",x"6d",x"49",x"24",x"6d",x"db",x"92",x"92",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"48",x"24",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"6d",x"db",x"b4",x"b4",x"92",x"92",x"b4",x"90",x"90",x"6d",x"49",x"24",x"49",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"49",x"48",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"90",x"90",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",
--x"6d",x"b4",x"b4",x"90",x"b6",x"92",x"90",x"6c",x"6c",x"6d",x"49",x"24",x"49",x"db",x"92",x"92",x"90",x"6d",x"92",x"6d",x"6d",x"49",x"48",x"24",x"25",x"49",x"6d",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"d4",x"d4",x"b4",x"90",x"b6",x"b6",x"d8",x"b4",x"b6",x"d4",x"b4",x"90",x"b6",x"6d",x"49",x"49",
--x"6d",x"b4",x"90",x"6d",x"92",x"92",x"92",x"6c",x"6c",x"6d",x"24",x"25",x"49",x"db",x"b6",x"92",x"90",x"6d",x"b6",x"92",x"6d",x"49",x"48",x"24",x"24",x"49",x"6c",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"90",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"b4",x"90",x"90",x"90",x"b6",x"b6",x"d8",x"b4",x"b6",x"b6",x"b4",x"b4",x"b4",x"90",x"6d",x"25",x"49",
--x"6d",x"b4",x"90",x"6d",x"b6",x"92",x"92",x"92",x"92",x"49",x"24",x"25",x"49",x"db",x"92",x"b6",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"48",x"24",x"24",x"49",x"6c",x"d4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"90",x"92",x"b6",x"92",x"b4",x"90",x"b6",x"92",x"d4",x"d4",x"b4",x"6d",x"92",x"b6",x"b4",x"90",x"b4",x"90",x"6d",x"49",x"25",x"49",
--x"6d",x"b4",x"90",x"92",x"92",x"b6",x"92",x"b6",x"92",x"49",x"24",x"49",x"49",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"6d",x"49",x"48",x"24",x"24",x"49",x"25",x"b4",x"b4",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"6c",x"92",x"b6",x"b6",x"b6",x"90",x"90",x"b6",x"b6",x"92",x"b6",x"92",x"b6",x"d4",x"b4",x"b4",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"b4",x"6d",x"6d",x"49",x"25",x"49",
--x"49",x"90",x"6d",x"92",x"b6",x"92",x"b6",x"92",x"6d",x"49",x"24",x"49",x"49",x"da",x"92",x"92",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"92",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"6c",x"6c",x"6d",x"b6",x"b6",x"b6",x"92",x"6d",x"92",x"b6",x"92",x"92",x"b6",x"d4",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"92",x"92",x"b4",x"6d",x"6d",x"49",x"25",x"49",
--x"49",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"25",x"49",x"49",x"b6",x"b6",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"b6",x"90",x"6c",x"6c",x"6c",x"6c",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"92",x"92",x"d4",x"d4",x"92",x"92",x"6d",x"6d",x"92",x"92",x"d8",x"b4",x"b6",x"b6",x"92",x"b4",x"6d",x"6d",x"49",x"25",x"49",
--x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"92",x"92",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"da",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"90",x"b6",x"b6",x"b6",x"92",x"b6",x"d4",x"b6",x"92",x"92",x"b6",x"92",x"92",x"92",x"b6",x"b4",x"90",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"49",
--x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"da",x"6d",x"6d",x"92",x"92",x"b4",x"b4",x"90",x"b6",x"92",x"92",x"b6",x"92",x"b6",x"b6",x"b6",x"92",x"b4",x"b6",x"b4",x"b6",x"92",x"b6",x"b4",x"90",x"92",x"b6",x"b6",x"92",x"b4",x"b4",x"6d",x"49",x"24",x"49",
--x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"25",x"92",x"da",x"b6",x"92",x"b6",x"92",x"b6",x"b4",x"b4",x"6c",x"92",x"b6",x"92",x"b6",x"92",x"92",x"92",x"d8",x"b4",x"6c",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"6d",x"49",x"24",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"90",x"6c",x"6c",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"d8",x"b4",x"6c",x"b6",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"92",x"92",x"d4",x"92",x"92",x"92",x"6d",x"49",x"24",x"49",
--x"49",x"6d",x"b6",x"d4",x"d4",x"d4",x"90",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"6d",x"6d",x"6d",x"92",x"b4",x"b6",x"6c",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"49",
--x"49",x"b6",x"d4",x"d8",x"d4",x"d4",x"d4",x"d4",x"b4",x"90",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",
--x"49",x"b6",x"d4",x"d8",x"b4",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b4",x"d8",x"d8",x"d4",x"d4",x"d4",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",
--x"49",x"b6",x"b6",x"92",x"b4",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",
--x"49",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"90",x"90",x"90",x"92",x"92",x"b6",x"db",x"d8",x"d8",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"d8",x"b4",x"90",x"b6",x"b6",x"da",x"b6",x"da",x"b6",x"b6",x"d4",x"90",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"92",x"d8",x"90",x"92",x"6d",x"6d",x"24",x"49",x"49",x"49",x"90",x"b4",x"b4",x"b4",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6c",x"b4",x"90",x"90",x"6c",x"6c",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
--x"49",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"b4",x"90",x"48",x"b6",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"b6",x"b6",x"da",x"b6",x"6d",x"b6",x"da",x"b6",x"92",x"92",x"6d",x"49",x"24",x"49",x"49",x"49",x"b4",x"90",x"90",x"90",x"6d",x"db",x"db",x"b6",x"49",x"49",x"90",x"d4",x"d4",x"d4",x"90",x"6d",x"d4",x"b6",x"b6",x"da",x"d4",x"b6",x"92",x"6d",x"49",x"49",x"49",
--x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"90",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"90",x"90",x"6c",x"6d",x"b6",x"b6",x"b6",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"92",x"d4",x"90",x"6d",x"b6",x"db",x"92",x"24",x"49",
--x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"b6",x"90",x"6c",x"6d",x"92",x"6d",x"92",x"92",x"6d",x"49",x"92",x"92",x"b6",x"92",x"b6",x"d4",x"d4",x"b6",x"b6",x"90",x"90",x"6d",x"92",x"b6",x"49",x"24",x"49",
--x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"48",x"48",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"b6",x"d4",x"d4",x"90",x"6d",x"b6",x"90",x"6d",x"6d",x"92",x"92",x"49",x"24",x"49",
--x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"48",x"48",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6c",x"48",x"49",x"49",x"49",x"6c",x"48",x"49",x"49",x"49",x"49",x"49",x"24",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",
--x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"
--
--);

constant ROM: rom_type := (


--00 BlueStone



x"383838",x"000070",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000070",x"383838",x"383838",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"000088",x"383838",x"383838",x"000070",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000070",x"2c2c2c",
x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"202020",x"202020",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"202020",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"202020",
x"000000",x"0000a4",x"0000a4",x"0000a4",x"000088",x"0000a4",x"00007c",x"0000a4",x"0000a4",x"000098",x"00007c",x"000098",x"000098",x"00007c",x"000098",x"000098",x"00007c",x"0000a4",x"00007c",x"000070",x"000070",x"000058",x"000000",x"202020",x"0000bc",x"0000a4",x"0000bc",x"0000b0",x"00007c",x"0000a4",x"0000bc",x"000098",x"000070",x"000070",x"000098",x"000088",x"0000a4",x"0000a4",x"000088",x"000070",x"000088",x"0000a4",x"0000bc",x"0000a4",x"000088",x"000098",x"0000a4",x"0000bc",x"0000bc",x"0000a4",x"000098",x"000070",x"000000",x"202020",x"0000b0",x"0000bc",x"0000a4",x"000098",x"0000a4",x"0000b0",x"0000b0",x"000098",x"00007c",x"000000",
x"000000",x"0000a4",x"000098",x"00007c",x"000088",x"000098",x"000098",x"000098",x"00007c",x"00007c",x"0000a4",x"000098",x"0000a4",x"000064",x"000098",x"000098",x"00007c",x"000070",x"00007c",x"00007c",x"000070",x"000064",x"000000",x"202020",x"0000bc",x"0000bc",x"0000a4",x"000098",x"000098",x"000098",x"000070",x"000098",x"000058",x"000070",x"000058",x"000058",x"00007c",x"0000a4",x"0000a4",x"000064",x"000070",x"000070",x"000064",x"000070",x"000070",x"000058",x"000070",x"000088",x"000088",x"000070",x"000064",x"000070",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"00007c",x"000098",x"0000a4",x"0000a4",x"000058",x"000000",
x"000000",x"0000a4",x"000088",x"0000a4",x"000070",x"0000c8",x"0000c8",x"000098",x"00007c",x"00007c",x"00007c",x"000098",x"000088",x"000088",x"00007c",x"000064",x"000058",x"00007c",x"000070",x"000058",x"000058",x"000064",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000b0",x"0000a4",x"0000b0",x"0000bc",x"0000bc",x"0000b0",x"0000a4",x"00007c",x"00007c",x"000000",
x"000000",x"0000a4",x"000088",x"00007c",x"0000a4",x"0000c8",x"0000c8",x"000064",x"00007c",x"00007c",x"00007c",x"0000a4",x"000098",x"000098",x"000098",x"000088",x"000070",x"000070",x"00007c",x"000058",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"0000b0",x"0000bc",x"0000a4",x"0000b0",x"0000a4",x"00007c",x"00007c",x"000064",x"000058",x"000000",
x"000000",x"0000a4",x"000098",x"000098",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"000098",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000098",x"000070",x"000070",x"000064",x"000058",x"000064",x"000070",x"000064",x"000000",x"202020",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000a4",x"000098",x"000098",x"0000bc",x"000098",x"000098",x"0000b0",x"000098",x"000098",x"0000b0",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000098",x"000064",x"202020",x"202020",x"0000b0",x"000098",x"000098",x"0000a4",x"00007c",x"000088",x"000088",x"000064",x"000064",x"000000",
x"000000",x"0000a4",x"0000a4",x"000098",x"0000a4",x"0000b0",x"0000b0",x"0000a4",x"000098",x"00007c",x"000064",x"0000a4",x"0000a4",x"000098",x"000088",x"000088",x"00007c",x"000064",x"000064",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000bc",x"0000e0",x"0000c8",x"0000b0",x"0000a4",x"0000bc",x"0000a4",x"000098",x"000098",x"000098",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"000098",x"0000a4",x"000000",x"202020",x"0000a4",x"000098",x"000098",x"000088",x"000098",x"00007c",x"000064",x"000000",x"202020",x"0000b0",x"000098",x"000098",x"0000a4",x"000070",x"000088",x"000088",x"000088",x"000064",x"000000",
x"000000",x"0000a4",x"000098",x"00007c",x"000098",x"0000a4",x"0000a4",x"000088",x"000098",x"00007c",x"000098",x"000070",x"000070",x"000088",x"000088",x"000088",x"000070",x"00007c",x"00007c",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000c8",x"0000bc",x"0000c8",x"000098",x"0000b0",x"0000a4",x"0000a4",x"0000bc",x"000098",x"000098",x"0000a4",x"00007c",x"0000a4",x"00007c",x"000098",x"0000a4",x"00007c",x"000000",x"202020",x"0000a4",x"000098",x"000098",x"000098",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"0000b0",x"0000bc",x"0000a4",x"000098",x"0000a4",x"0000a4",x"000088",x"000088",x"000040",x"000000",
x"000000",x"0000a4",x"000088",x"000088",x"000088",x"0000a4",x"00007c",x"00007c",x"00007c",x"0000a4",x"0000a4",x"000070",x"000058",x"000064",x"000064",x"000070",x"000064",x"00007c",x"00007c",x"00007c",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"000098",x"000098",x"000098",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000088",x"000064",x"00007c",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"000098",x"00007c",x"00007c",x"000058",x"000058",x"000000",x"202020",x"0000bc",x"00007c",x"00007c",x"000098",x"0000a4",x"0000a4",x"000098",x"000058",x"000040",x"000000",
x"000000",x"000098",x"00007c",x"000088",x"0000a4",x"000088",x"000088",x"000070",x"000098",x"0000a4",x"0000a4",x"000070",x"000070",x"000064",x"000058",x"000064",x"000064",x"000064",x"00007c",x"00007c",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000bc",x"0000b0",x"0000b0",x"0000b0",x"000098",x"000098",x"0000b0",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"000064",x"000064",x"000088",x"00007c",x"00007c",x"000064",x"000058",x"000000",x"202020",x"0000a4",x"0000a4",x"000098",x"00007c",x"0000a4",x"00007c",x"000058",x"000000",x"202020",x"0000bc",x"00007c",x"0000bc",x"0000a4",x"00007c",x"000098",x"000098",x"000058",x"000040",x"000000",
x"000000",x"000098",x"000088",x"000098",x"00007c",x"00007c",x"0000a4",x"000088",x"000064",x"00007c",x"000058",x"00007c",x"000064",x"000058",x"000064",x"00007c",x"000040",x"000058",x"000040",x"000040",x"000064",x"000040",x"000000",x"202020",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000bc",x"0000b0",x"0000b0",x"0000a4",x"000064",x"000064",x"000070",x"0000a4",x"000064",x"000064",x"000040",x"000000",x"202020",x"0000a4",x"00007c",x"000088",x"000098",x"00007c",x"000058",x"000058",x"000000",x"202020",x"0000bc",x"0000bc",x"00007c",x"00007c",x"000064",x"000064",x"00007c",x"00007c",x"000040",x"000000",
x"000000",x"000098",x"00007c",x"000098",x"00007c",x"000064",x"000088",x"000088",x"00007c",x"000064",x"00007c",x"000064",x"00007c",x"000064",x"000040",x"000070",x"000070",x"000040",x"000040",x"000040",x"000064",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000a4",x"0000a4",x"000098",x"0000bc",x"000098",x"000098",x"0000a4",x"0000b0",x"0000b0",x"0000a4",x"000098",x"000098",x"00007c",x"00007c",x"000058",x"000058",x"000064",x"000000",x"202020",x"0000a4",x"000088",x"000088",x"000088",x"000070",x"000070",x"000064",x"000000",x"202020",x"0000bc",x"00007c",x"000070",x"000064",x"00007c",x"000064",x"00007c",x"00007c",x"000040",x"000000",
x"000000",x"000098",x"000098",x"00007c",x"00007c",x"00007c",x"000070",x"000064",x"000058",x"000058",x"000064",x"00007c",x"000064",x"000070",x"000064",x"000040",x"000040",x"000070",x"000040",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000e0",x"0000c8",x"000088",x"000088",x"000098",x"000098",x"000088",x"00007c",x"00007c",x"00007c",x"000088",x"000098",x"000088",x"00007c",x"000064",x"000064",x"000040",x"000000",x"202020",x"0000a4",x"0000a4",x"000088",x"000088",x"000070",x"000070",x"000064",x"000000",x"202020",x"0000bc",x"00007c",x"00007c",x"000070",x"000058",x"000058",x"000058",x"000058",x"000040",x"000000",
x"000000",x"000098",x"00007c",x"000098",x"000064",x"000064",x"000070",x"000064",x"00007c",x"000064",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000a4",x"0000bc",x"0000c8",x"0000c8",x"000088",x"000088",x"000088",x"0000a4",x"0000a4",x"00007c",x"000088",x"000088",x"00007c",x"000088",x"000070",x"00007c",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"00007c",x"000098",x"0000a4",x"000058",x"000058",x"000058",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"000098",x"000088",x"000088",x"0000a4",x"0000a4",x"0000a4",x"000088",x"000088",x"000098",x"000064",x"000064",x"00007c",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"000098",x"0000a4",x"000058",x"000064",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",
x"0000a4",x"0000bc",x"0000b0",x"0000a4",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000000",x"0000b0",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"000098",x"000098",x"000000",x"0000a4",x"0000b0",x"000098",x"0000a4",x"000088",x"000098",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"000098",x"000098",x"00007c",x"00007c",x"000058",x"000058",x"000040",x"000040",x"000000",x"202020",x"000098",x"0000a4",x"000098",x"0000a4",x"000098",x"000070",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000000",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",
x"0000bc",x"0000b0",x"0000a4",x"000098",x"0000a4",x"0000bc",x"0000b0",x"0000a4",x"000088",x"0000a4",x"0000a4",x"00007c",x"0000a4",x"000098",x"00007c",x"000000",x"0000b0",x"0000b0",x"000098",x"0000bc",x"0000bc",x"00007c",x"0000bc",x"000000",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000bc",x"0000a4",x"000098",x"0000a4",x"0000a4",x"0000a4",x"000088",x"000064",x"000070",x"00007c",x"000040",x"000040",x"000064",x"000058",x"000040",x"000000",x"202020",x"000098",x"000098",x"00007c",x"000070",x"00007c",x"000070",x"000058",x"000000",x"202020",x"0000a4",x"0000b0",x"000088",x"00007c",x"000000",x"0000bc",x"0000bc",x"0000a4",x"0000b0",x"0000bc",
x"0000bc",x"0000b0",x"000098",x"000098",x"000088",x"0000a4",x"0000a4",x"000088",x"00007c",x"000098",x"000098",x"00007c",x"00007c",x"000098",x"000098",x"000000",x"0000b0",x"0000bc",x"0000bc",x"0000b0",x"000098",x"00007c",x"00007c",x"000000",x"0000a4",x"0000b0",x"000098",x"0000a4",x"0000bc",x"0000a4",x"000088",x"00007c",x"000088",x"000088",x"000064",x"00007c",x"00007c",x"000070",x"000040",x"000040",x"000064",x"000040",x"000040",x"000000",x"202020",x"000098",x"000098",x"000058",x"000058",x"000058",x"000064",x"000040",x"000000",x"202020",x"0000a4",x"0000b0",x"0000b0",x"00007c",x"000000",x"0000bc",x"0000a4",x"0000b0",x"0000b0",x"0000b0",
x"0000b0",x"0000a4",x"000098",x"0000b0",x"0000b0",x"000098",x"000098",x"00007c",x"00007c",x"00007c",x"000098",x"00007c",x"00007c",x"00007c",x"00007c",x"000000",x"0000b0",x"0000bc",x"0000b0",x"0000b0",x"000098",x"000098",x"000064",x"000000",x"0000a4",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"000088",x"0000a4",x"00007c",x"00007c",x"000064",x"000070",x"000070",x"000058",x"000058",x"000058",x"000064",x"000064",x"000058",x"000040",x"000000",x"202020",x"000098",x"00007c",x"000058",x"000064",x"000058",x"000058",x"000040",x"000000",x"202020",x"0000a4",x"000088",x"00007c",x"000058",x"000000",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000b0",
x"0000a4",x"000088",x"000098",x"0000b0",x"0000bc",x"0000b0",x"00007c",x"00007c",x"000098",x"000098",x"00007c",x"000098",x"000058",x"00007c",x"00007c",x"000000",x"0000b0",x"0000bc",x"000098",x"00007c",x"000098",x"000098",x"000064",x"000000",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000098",x"000098",x"000098",x"00007c",x"000064",x"000058",x"000064",x"000064",x"000058",x"000064",x"000064",x"000058",x"000040",x"000040",x"000040",x"000000",x"202020",x"000098",x"00007c",x"000064",x"000058",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000a4",x"000058",x"000064",x"000058",x"000000",x"0000bc",x"0000bc",x"0000b0",x"0000b0",x"0000b0",
x"0000a4",x"0000a4",x"000088",x"000098",x"0000b0",x"0000d4",x"00007c",x"000098",x"00007c",x"00007c",x"000064",x"000064",x"000070",x"00007c",x"00007c",x"000000",x"0000b0",x"000098",x"0000bc",x"00007c",x"00007c",x"00007c",x"000064",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"000098",
x"0000b0",x"000088",x"00007c",x"000088",x"000098",x"0000a4",x"000098",x"00007c",x"00007c",x"000098",x"000064",x"000070",x"00007c",x"000058",x"000058",x"000000",x"0000b0",x"000098",x"000098",x"000064",x"00007c",x"00007c",x"000058",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"202020",x"202020",x"0000bc",x"0000a4",x"0000a4",x"000098",x"000098",
x"0000b0",x"0000a4",x"000088",x"000098",x"00007c",x"000098",x"00007c",x"000098",x"000098",x"00007c",x"000070",x"00007c",x"000064",x"00007c",x"000058",x"000000",x"0000b0",x"0000bc",x"000098",x"000088",x"000064",x"000058",x"000064",x"000000",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"000098",x"0000a4",x"202020",x"202020",x"0000b0",x"0000c8",x"0000b0",x"0000c8",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000000",x"202020",x"0000bc",x"0000b0",x"000098",x"000098",x"000098",
x"0000b0",x"0000b0",x"000098",x"000088",x"0000b0",x"000098",x"000098",x"000098",x"000098",x"00007c",x"00007c",x"000070",x"000058",x"000058",x"000058",x"000000",x"0000a4",x"0000bc",x"00007c",x"000088",x"000088",x"000064",x"000058",x"000000",x"202020",x"0000b0",x"0000bc",x"0000b0",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000bc",x"0000a4",x"0000b0",x"0000a4",x"0000bc",x"0000b0",x"00007c",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"00007c",x"0000a4",x"000058",x"000000",x"202020",x"0000b0",x"0000c8",x"0000b0",x"0000c8",x"0000c8",x"0000a4",x"000098",x"000088",x"000000",x"202020",x"0000bc",x"0000bc",x"000098",x"000098",x"000098",
x"0000b0",x"0000a4",x"000088",x"00007c",x"000088",x"0000b0",x"0000b0",x"000064",x"00007c",x"000098",x"000088",x"000088",x"000070",x"000058",x"000064",x"000000",x"0000a4",x"00007c",x"000064",x"000070",x"000070",x"000058",x"000064",x"000000",x"202020",x"0000b0",x"0000bc",x"0000a4",x"0000b0",x"0000c8",x"0000e0",x"0000e0",x"0000bc",x"0000d4",x"0000e0",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"000058",x"000000",x"202020",x"0000b0",x"0000c8",x"0000c8",x"0000c8",x"0000c8",x"0000a4",x"000088",x"00007c",x"000000",x"202020",x"0000bc",x"0000b0",x"0000bc",x"0000a4",x"0000a4",
x"0000a4",x"000098",x"00007c",x"000088",x"0000a4",x"0000b0",x"0000b0",x"0000a4",x"000098",x"00007c",x"000088",x"000088",x"000070",x"000058",x"000064",x"000000",x"000098",x"00007c",x"000058",x"000058",x"000058",x"000058",x"000064",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"0000bc",x"0000d4",x"0000d4",x"0000e0",x"0000bc",x"0000e0",x"0000d4",x"0000d4",x"0000b0",x"00007c",x"0000a4",x"00007c",x"00007c",x"0000a4",x"00007c",x"00007c",x"0000a4",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"0000c8",x"0000a4",x"000088",x"0000a4",x"000064",x"000000",x"202020",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"0000a4",
x"0000b0",x"000098",x"0000b0",x"000098",x"000098",x"0000a4",x"0000b0",x"0000a4",x"000064",x"00007c",x"000070",x"000070",x"000070",x"000058",x"000058",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000b0",x"0000bc",x"0000bc",x"0000b0",x"0000b0",x"0000c8",x"0000c8",x"0000a4",x"0000a4",x"0000d4",x"0000d4",x"0000a4",x"0000a4",x"00007c",x"00007c",x"00007c",x"000070",x"0000a4",x"00007c",x"00007c",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000c8",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000088",x"000064",x"000000",x"202020",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000b0",
x"0000a4",x"000088",x"000088",x"0000a4",x"0000a4",x"000098",x"0000a4",x"0000a4",x"000064",x"000070",x"000058",x"000064",x"000058",x"000040",x"000040",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"0000b0",x"0000b0",x"0000bc",x"0000b0",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"000088",x"000088",x"00007c",x"00007c",x"000058",x"000058",x"000058",x"000064",x"000000",x"202020",x"0000b0",x"0000c8",x"0000c8",x"0000a4",x"0000a4",x"000088",x"00007c",x"000070",x"000000",x"202020",x"0000bc",x"0000a4",x"0000a4",x"0000bc",x"0000b0",
x"0000a4",x"000098",x"000088",x"0000a4",x"0000a4",x"0000a4",x"000098",x"00007c",x"000070",x"000064",x"000058",x"000064",x"000064",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"202020",x"202020",x"0000b0",x"0000a4",x"0000a4",x"0000bc",x"0000b0",x"000088",x"000088",x"0000a4",x"0000bc",x"0000b0",x"00007c",x"0000a4",x"0000a4",x"00007c",x"000088",x"000088",x"000088",x"000070",x"000070",x"000070",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000c8",x"0000c8",x"000098",x"000098",x"0000a4",x"0000a4",x"000058",x"000000",x"202020",x"0000bc",x"0000a4",x"0000a4",x"0000b0",x"0000b0",
x"000098",x"000088",x"000098",x"000088",x"0000a4",x"0000a4",x"00007c",x"000064",x"000064",x"000058",x"000058",x"000058",x"000064",x"000040",x"000064",x"000000",x"202020",x"0000b0",x"0000b0",x"000088",x"0000a4",x"000098",x"000088",x"000000",x"202020",x"0000b0",x"0000bc",x"0000b0",x"0000bc",x"0000b0",x"000088",x"000088",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"0000a4",x"0000a4",x"0000a4",x"000070",x"000088",x"000088",x"000058",x"000070",x"000070",x"000070",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000c8",x"000098",x"000098",x"000098",x"0000a4",x"000058",x"000000",x"202020",x"0000bc",x"0000bc",x"000098",x"000098",x"00007c",
x"000098",x"000088",x"000088",x"00007c",x"000088",x"000088",x"00007c",x"000064",x"000064",x"000070",x"00007c",x"00007c",x"000064",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000a4",x"0000a4",x"000098",x"000088",x"000098",x"000000",x"202020",x"0000b0",x"0000bc",x"0000bc",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"000098",x"0000a4",x"00007c",x"00007c",x"00007c",x"0000a4",x"0000a4",x"000070",x"000058",x"000064",x"000058",x"000064",x"000070",x"000070",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"000088",x"0000b0",x"0000a4",x"0000a4",x"000064",x"000000",x"202020",x"0000bc",x"000088",x"000088",x"000098",x"000098",
x"000098",x"000088",x"0000a4",x"000098",x"000070",x"00007c",x"00007c",x"000070",x"000064",x"000070",x"00007c",x"00007c",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000b0",x"0000a4",x"000098",x"000088",x"000070",x"000064",x"000000",x"202020",x"0000b0",x"0000bc",x"0000a4",x"00007c",x"0000a4",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"00007c",x"000070",x"00007c",x"000064",x"000070",x"000070",x"000070",x"000058",x"000040",x"000040",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000c8",x"000088",x"0000b0",x"0000b0",x"000098",x"000064",x"000000",x"202020",x"0000bc",x"000088",x"000088",x"00007c",x"00007c",
x"000098",x"0000a4",x"000098",x"000088",x"000088",x"00007c",x"000064",x"000064",x"000058",x"00004c",x"00004c",x"000070",x"000064",x"000058",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"000088",x"0000b0",x"000088",x"000058",x"000000",x"202020",x"0000b0",x"0000a4",x"0000a4",x"0000bc",x"00007c",x"0000a4",x"0000a4",x"000098",x"00007c",x"000070",x"00007c",x"00007c",x"000064",x"000064",x"000070",x"000070",x"000064",x"000040",x"000040",x"000064",x"000064",x"000040",x"000000",x"202020",x"0000b0",x"0000a4",x"0000c8",x"0000a4",x"000088",x"000098",x"000098",x"000058",x"000000",x"202020",x"0000bc",x"0000bc",x"00007c",x"00007c",x"00007c",
x"00007c",x"000098",x"000098",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"000058",x"00004c",x"00004c",x"000058",x"000058",x"000064",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000b0",x"000070",x"000070",x"000064",x"000000",x"202020",x"0000b0",x"00007c",x"0000bc",x"00007c",x"0000a4",x"0000a4",x"00007c",x"00007c",x"000070",x"000064",x"00007c",x"00007c",x"00007c",x"000064",x"000064",x"000058",x"000058",x"000064",x"000064",x"000064",x"00004c",x"000040",x"000000",x"202020",x"0000b0",x"0000c8",x"0000a4",x"0000a4",x"000098",x"000058",x"000070",x"000064",x"000000",x"202020",x"0000bc",x"0000a4",x"0000a4",x"000098",x"000098",
x"00007c",x"000088",x"000088",x"00007c",x"000070",x"00007c",x"00007c",x"00007c",x"000058",x"000058",x"000064",x"000058",x"000058",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000a4",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000a4",x"0000bc",x"00007c",x"0000a4",x"0000a4",x"000070",x"000064",x"000064",x"000058",x"00007c",x"00007c",x"00007c",x"000064",x"000058",x"000058",x"000058",x"000058",x"00004c",x"00004c",x"00004c",x"000040",x"000000",x"202020",x"0000b0",x"0000c8",x"0000a4",x"000098",x"00007c",x"000098",x"000070",x"000058",x"000000",x"202020",x"0000bc",x"0000a4",x"0000a4",x"000098",x"000088",
x"00007c",x"000088",x"000064",x"000070",x"00007c",x"000064",x"00007c",x"00007c",x"000058",x"000064",x"000058",x"000040",x"000058",x"000064",x"000058",x"000000",x"202020",x"0000b0",x"000098",x"000098",x"000058",x"000088",x"000064",x"000000",x"202020",x"0000b0",x"0000a4",x"00007c",x"0000a4",x"0000a4",x"00007c",x"000058",x"000058",x"000058",x"000058",x"000064",x"000064",x"000064",x"000064",x"000058",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000c8",x"0000a4",x"00007c",x"000098",x"000098",x"00007c",x"000064",x"000000",x"202020",x"0000bc",x"000098",x"0000a4",x"0000a4",x"00007c",
x"00007c",x"000098",x"00007c",x"000064",x"00007c",x"000064",x"000070",x"000058",x"000064",x"000040",x"000040",x"000058",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"000098",x"000098",x"0000b0",x"000058",x"000064",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000a4",x"0000b0",x"0000a4",x"00007c",x"000064",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"0000bc",x"000098",x"000088",x"000088",x"00007c",
x"00007c",x"000088",x"000098",x"000088",x"000070",x"00007c",x"000070",x"000058",x"000058",x"000058",x"000040",x"000064",x"000040",x"000058",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"000088",x"0000b0",x"000088",x"000058",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"0000a4",x"0000b0",x"0000b0",x"0000a4",x"00007c",x"000058",x"000064",x"000040",x"000000",x"202020",x"0000bc",x"0000bc",x"000088",x"000088",x"00007c",
x"00007c",x"000098",x"000088",x"00007c",x"000064",x"000070",x"00007c",x"000070",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"000088",x"000088",x"000058",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"202020",x"202020",x"0000a4",x"0000b0",x"0000a4",x"0000bc",x"0000a4",x"00007c",x"000064",x"000040",x"000000",x"202020",x"0000bc",x"000098",x"000098",x"00007c",x"000088",
x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000b0",x"0000b0",x"00007c",x"00007c",x"000058",x"000058",x"000000",x"202020",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000088",x"00007c",x"0000bc",x"000098",x"0000a4",x"00007c",x"000000",x"202020",x"0000a4",x"0000c8",x"0000a4",x"0000a4",x"0000bc",x"000088",x"000058",x"000040",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",
x"202020",x"202020",x"202020",x"202020",x"202020",x"000058",x"000058",x"000070",x"000070",x"000088",x"000088",x"000088",x"00007c",x"000070",x"000064",x"202020",x"202020",x"0000a4",x"0000b0",x"00007c",x"00007c",x"00007c",x"000058",x"000000",x"202020",x"0000b0",x"0000bc",x"0000c8",x"0000c8",x"0000bc",x"0000a4",x"0000a4",x"0000b0",x"0000b0",x"0000c8",x"0000bc",x"000098",x"000098",x"0000a4",x"0000a4",x"000098",x"00007c",x"000088",x"00007c",x"000088",x"000098",x"00007c",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"000088",x"000088",x"000058",x"000040",x"000000",x"202020",x"000088",x"000098",x"000088",x"000088",x"000000",
x"202020",x"000098",x"0000a4",x"0000b0",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"202020",x"202020",x"0000a4",x"0000a4",x"000088",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"0000b0",x"0000bc",x"0000c8",x"0000c8",x"0000c8",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000bc",x"0000bc",x"00007c",x"00007c",x"00007c",x"00007c",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000098",x"00007c",x"000064",x"000000",x"202020",x"0000a4",x"0000c8",x"0000a4",x"00007c",x"000070",x"000058",x"000058",x"000040",x"000000",x"202020",x"000098",x"000098",x"00007c",x"00007c",x"000000",
x"202020",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000a4",x"0000b0",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"0000bc",x"000000",x"202020",x"0000a4",x"0000a4",x"000098",x"000058",x"000064",x"000064",x"000000",x"202020",x"0000b0",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000d4",x"0000d4",x"0000b0",x"0000b0",x"0000b0",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000098",x"00007c",x"00007c",x"000070",x"000098",x"000064",x"000000",x"202020",x"0000a4",x"0000b0",x"000088",x"000070",x"000064",x"000058",x"000070",x"000040",x"000000",x"202020",x"000098",x"00007c",x"000070",x"000070",x"000000",
x"202020",x"0000a4",x"0000bc",x"0000b0",x"0000b0",x"0000d4",x"0000d4",x"0000b0",x"0000bc",x"0000bc",x"0000bc",x"000098",x"0000a4",x"0000bc",x"0000bc",x"000000",x"202020",x"0000a4",x"000098",x"000088",x"000058",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000bc",x"0000bc",x"0000b0",x"0000bc",x"0000d4",x"0000d4",x"0000d4",x"00007c",x"0000a4",x"000098",x"00007c",x"00007c",x"000070",x"000070",x"000070",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"000070",x"000064",x"000070",x"000058",x"000058",x"000040",x"000000",x"202020",x"000098",x"000070",x"00007c",x"000058",x"000000",
x"202020",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"0000d4",x"0000d4",x"0000bc",x"000098",x"000098",x"0000a4",x"0000bc",x"0000bc",x"000098",x"0000b0",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"0000a4",x"0000b0",x"0000bc",x"0000b0",x"0000bc",x"0000bc",x"0000d4",x"0000d4",x"0000bc",x"0000a4",x"0000a4",x"000098",x"00007c",x"000070",x"000070",x"000064",x"000064",x"000058",x"00007c",x"00007c",x"00007c",x"000064",x"000000",x"202020",x"000088",x"00007c",x"00007c",x"000058",x"000058",x"000058",x"000064",x"000040",x"000000",x"202020",x"000088",x"00007c",x"000070",x"000058",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000b0",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"000098",x"000098",x"000098",x"0000bc",x"0000a4",x"000088",x"000088",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"0000a4",x"0000a4",x"0000b0",x"0000c8",x"000098",x"000098",x"0000bc",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"00007c",x"000064",x"000064",x"00007c",x"000064",x"000058",x"00004c",x"00004c",x"000000",x"202020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"202020",x"000088",x"000070",x"000058",x"000064",x"000000",
x"202020",x"0000bc",x"0000bc",x"0000b0",x"000098",x"000088",x"0000b0",x"0000b0",x"0000a4",x"000098",x"000098",x"0000a4",x"0000bc",x"0000bc",x"0000a4",x"000000",x"202020",x"0000bc",x"0000bc",x"0000b0",x"0000a4",x"0000a4",x"000098",x"202020",x"202020",x"0000a4",x"0000a4",x"0000c8",x"0000c8",x"000098",x"000098",x"000098",x"0000b0",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"00007c",x"000098",x"000088",x"000070",x"000064",x"000064",x"000058",x"000058",x"000040",x"000040",x"000000",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"000000",
x"202020",x"0000bc",x"0000bc",x"000098",x"0000a4",x"0000bc",x"0000b0",x"000088",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"00007c",x"0000a4",x"0000a4",x"000000",x"202020",x"0000bc",x"00007c",x"0000bc",x"000088",x"000098",x"000088",x"000000",x"202020",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000b0",x"000098",x"000098",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"00007c",x"00007c",x"00007c",x"00007c",x"000064",x"000064",x"000064",x"000058",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"000000",
x"202020",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"000088",x"0000bc",x"000088",x"0000b0",x"00007c",x"00007c",x"0000a4",x"000088",x"0000a4",x"000000",x"202020",x"0000bc",x"0000a4",x"0000b0",x"0000b0",x"000098",x"00007c",x"000000",x"202020",x"0000a4",x"0000b0",x"0000a4",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"00007c",x"000088",x"000070",x"000058",x"000064",x"000064",x"000064",x"000070",x"000058",x"00004c",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"0000b0",x"0000a4",x"000088",x"0000bc",x"0000a4",x"0000a4",x"00007c",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000bc",x"000098",x"0000a4",x"0000a4",x"0000bc",x"0000b0",x"000098",x"00007c",x"00004c",x"00007c",x"0000a4",x"0000a4",x"000000",x"202020",x"0000bc",x"0000bc",x"00007c",x"0000a4",x"00007c",x"000070",x"000000",x"202020",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"000098",x"0000a4",x"0000bc",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"000058",x"000058",x"000058",x"000058",x"000064",x"000070",x"000070",x"000064",x"000000",x"202020",x"0000b0",x"0000a4",x"0000b0",x"0000d4",x"0000d4",x"0000b0",x"0000b0",x"0000b0",x"000098",x"0000a4",x"0000a4",x"0000a4",x"000098",x"00007c",x"000000",
x"202020",x"0000bc",x"0000b0",x"000098",x"000098",x"0000bc",x"0000e0",x"0000bc",x"0000a4",x"000088",x"0000a4",x"00007c",x"00007c",x"0000a4",x"0000a4",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"0000a4",x"00007c",x"0000a4",x"000000",x"202020",x"0000a4",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"0000bc",x"000088",x"000088",x"0000bc",x"0000bc",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"000070",x"000058",x"000058",x"000064",x"000058",x"00004c",x"00004c",x"00004c",x"000000",x"202020",x"0000b0",x"0000bc",x"0000bc",x"0000d4",x"0000c8",x"0000c8",x"0000b0",x"0000b0",x"000088",x"000088",x"0000a4",x"000098",x"00007c",x"000064",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000bc",x"0000a4",x"0000e0",x"4040fc",x"0000e0",x"000098",x"000098",x"0000a4",x"000098",x"000088",x"00007c",x"000088",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"00007c",x"0000a4",x"000070",x"000000",x"202020",x"0000a4",x"0000a4",x"0000bc",x"000098",x"000098",x"00007c",x"00007c",x"00007c",x"000088",x"0000a4",x"0000a4",x"0000a4",x"00007c",x"00007c",x"00007c",x"000064",x"000064",x"000058",x"000058",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"000098",x"0000bc",x"000098",x"0000c8",x"0000c8",x"0000b0",x"0000b0",x"0000a4",x"0000a4",x"00007c",x"00007c",x"00007c",x"000058",x"000000",
x"202020",x"0000bc",x"0000b0",x"0000bc",x"0000b0",x"0000bc",x"0000e0",x"0000bc",x"0000a4",x"00007c",x"0000a4",x"0000a4",x"00004c",x"00004c",x"000064",x"000000",x"202020",x"0000bc",x"0000a4",x"0000b0",x"0000b0",x"00007c",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"0000bc",x"0000a4",x"000088",x"000088",x"00007c",x"00007c",x"00007c",x"000088",x"00007c",x"000088",x"000058",x"000058",x"000098",x"000098",x"000070",x"000070",x"000058",x"00004c",x"000040",x"000040",x"000000",x"202020",x"0000b0",x"0000bc",x"0000b0",x"000098",x"000098",x"000098",x"0000a4",x"0000a4",x"00007c",x"00007c",x"00007c",x"00007c",x"000058",x"000064",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000bc",x"0000b0",x"0000b0",x"0000b0",x"000088",x"000088",x"000088",x"00007c",x"000070",x"00004c",x"00004c",x"000064",x"000000",x"202020",x"0000bc",x"0000bc",x"0000b0",x"000098",x"000088",x"000064",x"000000",x"202020",x"0000a4",x"000098",x"0000bc",x"0000bc",x"000098",x"0000bc",x"00007c",x"00007c",x"000088",x"00007c",x"00007c",x"000088",x"00007c",x"000058",x"000098",x"000098",x"000088",x"000070",x"000070",x"000064",x"000058",x"000064",x"000000",x"202020",x"0000b0",x"0000b0",x"0000a4",x"000098",x"000098",x"000098",x"0000a4",x"00007c",x"000070",x"000064",x"00007c",x"000058",x"000058",x"000064",x"000000",
x"202020",x"0000a4",x"0000bc",x"0000b0",x"0000b0",x"0000a4",x"00007c",x"00007c",x"000098",x"0000a4",x"000098",x"000098",x"00007c",x"000064",x"000064",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"000088",x"000088",x"00007c",x"000000",x"202020",x"0000a4",x"0000bc",x"000098",x"0000a4",x"0000bc",x"0000a4",x"000088",x"00007c",x"000070",x"000070",x"000088",x"000088",x"000058",x"000058",x"00007c",x"000098",x"000098",x"00007c",x"000070",x"000058",x"000058",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"000098",x"0000a4",x"000098",x"000098",x"0000a4",x"00007c",x"000070",x"000064",x"000070",x"00007c",x"000058",x"000058",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000bc",x"0000b0",x"000088",x"000088",x"0000b0",x"00007c",x"0000a4",x"0000a4",x"000098",x"000070",x"00007c",x"000058",x"000000",x"202020",x"0000bc",x"0000a4",x"0000bc",x"00007c",x"00007c",x"00007c",x"000000",x"202020",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000088",x"0000a4",x"0000a4",x"000070",x"000070",x"000058",x"000070",x"000058",x"000058",x"00007c",x"00007c",x"00007c",x"000064",x"000058",x"000058",x"000040",x"000000",x"202020",x"0000b0",x"0000b0",x"0000bc",x"0000b0",x"000088",x"0000b0",x"0000b0",x"000098",x"00007c",x"000064",x"000098",x"000098",x"000058",x"000040",x"000000",
x"202020",x"0000bc",x"0000a4",x"0000bc",x"0000a4",x"000098",x"000088",x"00007c",x"000064",x"000088",x"0000a4",x"0000a4",x"000098",x"000070",x"000064",x"000000",x"202020",x"0000bc",x"0000bc",x"0000a4",x"000064",x"000064",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"0000a4",x"000098",x"000098",x"00007c",x"000088",x"0000a4",x"0000a4",x"0000a4",x"000070",x"000064",x"000070",x"000070",x"000058",x"00004c",x"00004c",x"00004c",x"000064",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000bc",x"0000bc",x"0000b0",x"000088",x"0000a4",x"0000b0",x"0000b0",x"0000b0",x"000098",x"00007c",x"000098",x"000098",x"00007c",x"000040",x"000000",
x"202020",x"0000b0",x"0000a4",x"000088",x"000088",x"000088",x"0000a4",x"000064",x"00004c",x"000064",x"000088",x"000098",x"000098",x"000070",x"000070",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"00007c",x"000070",x"000058",x"000000",x"202020",x"0000a4",x"0000b0",x"0000a4",x"000098",x"000098",x"0000bc",x"0000a4",x"00007c",x"0000a4",x"0000a4",x"000058",x"000058",x"000070",x"000070",x"000064",x"000058",x"000040",x"000040",x"000058",x"000040",x"000040",x"000040",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"000088",x"0000a4",x"0000a4",x"0000b0",x"0000b0",x"000098",x"00007c",x"00007c",x"00007c",x"00007c",x"000040",x"000000",
x"202020",x"0000b0",x"0000a4",x"000070",x"000064",x"000088",x"000064",x"0000a4",x"00007c",x"00007c",x"000098",x"000058",x"000064",x"000058",x"000058",x"000000",x"202020",x"0000b0",x"0000a4",x"000064",x"000064",x"000064",x"000058",x"000000",x"202020",x"0000a4",x"0000b0",x"0000bc",x"00007c",x"0000bc",x"0000bc",x"0000a4",x"000058",x"000064",x"000064",x"000064",x"000058",x"000058",x"00004c",x"00004c",x"00004c",x"000040",x"000040",x"00004c",x"000058",x"000040",x"000040",x"000000",x"202020",x"0000bc",x"0000b0",x"0000a4",x"0000bc",x"0000a4",x"0000a4",x"00007c",x"000088",x"000070",x"000070",x"00007c",x"00007c",x"000058",x"000040",x"000000",
x"202020",x"0000a4",x"0000a4",x"000088",x"000088",x"000064",x"000088",x"000058",x"000064",x"000058",x"000064",x"000070",x"000064",x"000070",x"000064",x"000000",x"202020",x"0000b0",x"0000a4",x"000088",x"000070",x"000064",x"000064",x"000000",x"202020",x"0000a4",x"0000a4",x"0000b0",x"0000bc",x"0000a4",x"00007c",x"000098",x"000058",x"000064",x"000064",x"000064",x"000058",x"000058",x"000040",x"000040",x"000070",x"000070",x"000064",x"000040",x"00004c",x"000040",x"000058",x"000000",x"202020",x"0000bc",x"0000bc",x"0000bc",x"000098",x"0000a4",x"00007c",x"00007c",x"000070",x"00007c",x"00007c",x"000070",x"000064",x"000040",x"000064",x"000000",
x"202020",x"0000a4",x"000098",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000070",x"000070",x"000070",x"000070",x"00007c",x"00007c",x"00007c",x"202020",x"202020",x"0000a4",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"202020",x"202020",x"0000a4",x"0000a4",x"000098",x"0000a4",x"000098",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000070",x"000064",x"000058",x"000058",x"00007c",x"00007c",x"00007c",x"00007c",x"000058",x"000058",x"000070",x"202020",x"202020",x"0000bc",x"0000a4",x"0000a4",x"00007c",x"000098",x"0000a4",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"000070",x"000070",x"00007c",x"000000",
x"383838",x"000088",x"000088",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"383838",x"383838",x"000088",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"383838",x"383838",x"0000a4",x"0000c8",x"000088",x"000088",x"000088",x"000088",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"383838",x"383838",x"0000bc",x"000088",x"000088",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"00007c",x"202020",
x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"383838",


--01 Eagle



x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",
x"545454",x"383838",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"484848",x"383838",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"484848",x"484848",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"383838",
x"383838",x"ec0000",x"ec0000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"a40000",x"484848",x"484848",x"545454",x"ec0000",x"ec0000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"a40000",x"484848",x"383838",x"545454",x"ec0000",x"ec0000",x"ec0000",x"ec0000",x"e00000",x"e00000",x"e00000",x"e00000",x"e00000",x"e00000",x"d40000",x"d40000",x"d40000",x"d40000",x"d40000",x"c80000",x"c80000",x"c80000",x"c80000",x"bc0000",x"bc0000",x"bc0000",x"a40000",x"484848",
x"484848",x"fcf400",x"c80000",x"b00000",x"b00000",x"d40000",x"880000",x"a40000",x"d40000",x"880000",x"c80000",x"a40000",x"640000",x"2c2c2c",x"484848",x"545454",x"ec0000",x"bc0000",x"880000",x"bc0000",x"880000",x"bc0000",x"880000",x"bc0000",x"7c0000",x"bc0000",x"980000",x"bc0000",x"980000",x"bc0000",x"7c0000",x"bc0000",x"7c0000",x"bc0000",x"c80000",x"a40000",x"700000",x"2c2c2c",x"484848",x"383838",x"d40000",x"a40000",x"c80000",x"b00000",x"c80000",x"b00000",x"b00000",x"c80000",x"700000",x"c80000",x"7c0000",x"c80000",x"b00000",x"c80000",x"880000",x"b00000",x"a40000",x"7c0000",x"c80000",x"980000",x"c80000",x"a40000",x"fcf400",x"2c2c2c",
x"e4d800",x"ccc400",x"848400",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"ccc400",x"ccc400",x"706c00",
x"a86840",x"9c9c00",x"585400",x"707070",x"707070",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"707070",x"707070",x"707070",x"706c00",x"e88c58",x"585400",
x"484848",x"543c1c",x"a40000",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"7c7c7c",x"707070",x"7c7c7c",x"7c7c7c",x"580000",x"a86840",x"2c2c2c",
x"484848",x"bc0000",x"7c0000",x"989898",x"7c7c7c",x"fc2020",x"a40000",x"400000",x"400000",x"545454",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"700000",x"a40000",x"b00000",x"fc0000",x"e00000",x"7c7c7c",x"400000",x"400000",x"400000",x"7c7c7c",x"c0c0c0",x"707070",x"580000",x"400000",x"2c2c2c",
x"484848",x"bc0000",x"a40000",x"a8a8a8",x"7c7c7c",x"a40000",x"c0c0c0",x"989898",x"707070",x"400000",x"7c7c7c",x"a8a8a8",x"c0c0c0",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"7c7c7c",x"400000",x"7c7c7c",x"707070",x"989898",x"fc2020",x"7c7c7c",x"707070",x"580000",x"400000",x"2c2c2c",
x"484848",x"7c0000",x"640000",x"b4b4b4",x"989898",x"400000",x"989898",x"c0c0c0",x"989898",x"7c7c7c",x"8c8c8c",x"989898",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"a8a8a8",x"d0d0d0",x"c0c0c0",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"6c0070",x"646464",x"c0c0c0",x"b4b4b4",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"707070",x"a8a8a8",x"d0d0d0",x"a40000",x"707070",x"7c7c7c",x"400000",x"400000",x"2c2c2c",
x"484848",x"484848",x"2c2c2c",x"d0d0d0",x"a8a8a8",x"400000",x"989898",x"a8a8a8",x"c0c0c0",x"989898",x"7c7c7c",x"7c7c7c",x"989898",x"989898",x"545454",x"580058",x"707070",x"a8a8a8",x"d0d0d0",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"8c8c8c",x"646464",x"600064",x"500050",x"989898",x"a8a8a8",x"a8a8a8",x"989898",x"989898",x"a8a8a8",x"d0d0d0",x"7c7c7c",x"400000",x"7c7c7c",x"989898",x"202020",x"202020",x"2c2c2c",
x"545454",x"383838",x"383838",x"d0d0d0",x"b4b4b4",x"545454",x"707070",x"989898",x"b4b4b4",x"c0c0c0",x"989898",x"7c7c7c",x"7c7c7c",x"8c8c8c",x"500050",x"580058",x"580058",x"580058",x"7c7c7c",x"a8a8a8",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"b4b4b4",x"500050",x"707070",x"545454",x"500050",x"500050",x"500050",x"500050",x"b45400",x"cc6000",x"fc7800",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"8c8c8c",x"646464",x"600064",x"580058",x"500050",x"500050",x"989898",x"989898",x"989898",x"989898",x"a8a8a8",x"d0d0d0",x"c0c0c0",x"646464",x"545454",x"8c8c8c",x"a8a8a8",x"202020",x"2c2c2c",x"2c2c2c",
x"ec0000",x"d40000",x"d40000",x"b4b4b4",x"d0d0d0",x"400000",x"7c7c7c",x"989898",x"a8a8a8",x"b4b4b4",x"c0c0c0",x"989898",x"707070",x"646464",x"484848",x"480048",x"500050",x"500050",x"580058",x"580058",x"7c7c7c",x"a8a8a8",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"500050",x"b45400",x"b45400",x"cc6000",x"fc8820",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"646464",x"600064",x"580058",x"500050",x"500050",x"500050",x"484848",x"989898",x"989898",x"989898",x"a8a8a8",x"c0c0c0",x"c0c0c0",x"a8a8a8",x"7c7c7c",x"400000",x"989898",x"a8a8a8",x"580000",x"580000",x"d40000",
x"b00000",x"880000",x"880000",x"b4b4b4",x"d0d0d0",x"700000",x"989898",x"8c8c8c",x"989898",x"a8a8a8",x"b4b4b4",x"646464",x"580058",x"707070",x"646464",x"484848",x"480048",x"480048",x"500050",x"500050",x"580058",x"580058",x"580058",x"7c7c7c",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b45400",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"646464",x"600064",x"600064",x"580058",x"580058",x"500050",x"500050",x"500050",x"484848",x"707070",x"707070",x"500050",x"646464",x"a8a8a8",x"c0c0c0",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"400000",x"a8a8a8",x"b4b4b4",x"580000",x"580000",x"b00000",
x"880000",x"a40000",x"880000",x"b4b4b4",x"d0d0d0",x"b00000",x"a8a8a8",x"989898",x"8c8c8c",x"989898",x"646464",x"6c0070",x"600064",x"484848",x"707070",x"646464",x"484848",x"480048",x"480048",x"480048",x"480048",x"840084",x"580058",x"580058",x"580058",x"707070",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"8c8c8c",x"b4b4b4",x"8c8c8c",x"646464",x"600064",x"600064",x"580058",x"840084",x"500050",x"500050",x"500050",x"480048",x"484848",x"707070",x"545454",x"6c0070",x"600064",x"600064",x"646464",x"a8a8a8",x"989898",x"7c7c7c",x"8c8c8c",x"700000",x"a8a8a8",x"b4b4b4",x"580000",x"580000",x"980000",
x"700000",x"a40000",x"a40000",x"b4b4b4",x"b4b4b4",x"980000",x"b4b4b4",x"989898",x"8c8c8c",x"8c8c8c",x"480048",x"600064",x"6c0070",x"600064",x"580058",x"484848",x"646464",x"484848",x"383838",x"480048",x"480048",x"6c0070",x"480048",x"580058",x"580058",x"580058",x"580058",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"580058",x"600064",x"600064",x"580058",x"500050",x"6c0070",x"480048",x"480048",x"383838",x"484848",x"646464",x"484848",x"500050",x"600064",x"600064",x"6c0070",x"6c0070",x"989898",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"700000",x"a8a8a8",x"b4b4b4",x"580000",x"580000",x"7c0000",
x"a40000",x"880000",x"880000",x"b4b4b4",x"b4b4b4",x"880000",x"c0c0c0",x"a8a8a8",x"989898",x"8c8c8c",x"480048",x"480048",x"600064",x"6c0070",x"600064",x"600064",x"580058",x"484848",x"545454",x"383838",x"400040",x"400040",x"480048",x"480048",x"480048",x"580058",x"545454",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"545454",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"383838",x"484848",x"484848",x"480048",x"500050",x"580058",x"600064",x"6c0070",x"6c0070",x"6c0070",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"700000",x"a8a8a8",x"b4b4b4",x"580000",x"580000",x"7c0000",
x"700000",x"a40000",x"640000",x"b4b4b4",x"b4b4b4",x"700000",x"d0d0d0",x"b4b4b4",x"a8a8a8",x"989898",x"484848",x"480048",x"480048",x"600064",x"6c0070",x"6c0070",x"600064",x"580058",x"480048",x"400040",x"400040",x"400040",x"400040",x"480048",x"480048",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"480048",x"480048",x"480048",x"400040",x"400040",x"400040",x"480048",x"480048",x"500050",x"580058",x"600064",x"6c0070",x"6c0070",x"6c0070",x"545454",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"989898",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"880000",
x"700000",x"b00000",x"640000",x"b4b4b4",x"b4b4b4",x"700000",x"d0d0d0",x"c0c0c0",x"b4b4b4",x"989898",x"646464",x"484848",x"480048",x"580058",x"600064",x"600064",x"6c0070",x"600064",x"580058",x"6c0070",x"400040",x"400040",x"400040",x"480048",x"8c8c8c",x"500050",x"707070",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"707070",x"480048",x"8c8c8c",x"480048",x"400040",x"400040",x"480048",x"580058",x"480048",x"480048",x"580058",x"600064",x"6c0070",x"6c0070",x"6c0070",x"545454",x"7c7c7c",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"700000",
x"400000",x"4c0000",x"4c0000",x"b4b4b4",x"b4b4b4",x"700000",x"d0d0d0",x"d0d0d0",x"646464",x"500050",x"707070",x"545454",x"545454",x"484848",x"580058",x"600064",x"600064",x"6c0070",x"580058",x"840084",x"500050",x"400040",x"400040",x"480048",x"500050",x"480048",x"500050",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"580058",x"6c0070",x"500050",x"580058",x"600064",x"600064",x"6c0070",x"545454",x"7c7c7c",x"646464",x"484848",x"484848",x"646464",x"989898",x"a8a8a8",x"700000",x"b4b4b4",x"b4b4b4",x"400000",x"580000",x"400000",
x"2c2c2c",x"2c2c2c",x"2c2c2c",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"d0d0d0",x"580058",x"500050",x"480048",x"484848",x"545454",x"545454",x"545454",x"484848",x"600064",x"600064",x"6c0070",x"580058",x"840084",x"500050",x"500050",x"500050",x"480048",x"500050",x"480048",x"7c7c7c",x"646464",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"646464",x"7c7c7c",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"6c0070",x"580058",x"580058",x"600064",x"600064",x"545454",x"8c8c8c",x"7c7c7c",x"646464",x"484848",x"400040",x"400040",x"480048",x"989898",x"a8a8a8",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"202020",x"2c2c2c",
x"545454",x"545454",x"484848",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"d0d0d0",x"600064",x"580058",x"500050",x"480048",x"480048",x"400040",x"383838",x"484848",x"484848",x"545454",x"646464",x"580058",x"580058",x"580058",x"580058",x"480048",x"480048",x"480048",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"500050",x"500050",x"580058",x"545454",x"646464",x"8c8c8c",x"7c7c7c",x"545454",x"500050",x"480048",x"400040",x"400040",x"400040",x"480048",x"a8a8a8",x"a8a8a8",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"2c2c2c",x"2c2c2c",
x"545454",x"ec0000",x"ec0000",x"c0c0c0",x"c0c0c0",x"7c0000",x"c0c0c0",x"b4b4b4",x"600064",x"600064",x"500050",x"500050",x"480048",x"400040",x"400040",x"400040",x"480048",x"480048",x"580058",x"9c009c",x"580058",x"580058",x"580058",x"480048",x"480048",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"480048",x"480048",x"480048",x"480048",x"480048",x"500050",x"580058",x"580058",x"9c009c",x"580058",x"580058",x"580058",x"500050",x"500050",x"480048",x"400040",x"400040",x"400040",x"400040",x"580058",x"a8a8a8",x"a8a8a8",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"2c2c2c",
x"545454",x"ec0000",x"880000",x"d0d0d0",x"d0d0d0",x"980000",x"d0d0d0",x"c0c0c0",x"580058",x"600064",x"580058",x"500050",x"480048",x"480048",x"400040",x"400040",x"400040",x"480048",x"480048",x"840084",x"580058",x"580058",x"580058",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"480048",x"480048",x"500050",x"500050",x"580058",x"580058",x"580058",x"9c009c",x"580058",x"580058",x"580058",x"500050",x"480048",x"480048",x"400040",x"400040",x"400040",x"480048",x"580058",x"989898",x"a8a8a8",x"7c0000",x"b4b4b4",x"b4b4b4",x"580000",x"400000",x"2c2c2c",
x"383838",x"ec0000",x"b00000",x"c0c0c0",x"c0c0c0",x"880000",x"c0c0c0",x"989898",x"707070",x"580058",x"600064",x"500050",x"500050",x"480048",x"400040",x"400040",x"480048",x"400040",x"480048",x"6c0070",x"580058",x"580058",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"545454",x"646464",x"707070",x"707070",x"646464",x"545454",x"545454",x"500050",x"500050",x"500050",x"580058",x"580058",x"580058",x"580058",x"580058",x"840084",x"580058",x"580058",x"500050",x"480048",x"480048",x"400040",x"400040",x"400040",x"400040",x"480048",x"707070",x"989898",x"a8a8a8",x"7c0000",x"b4b4b4",x"b4b4b4",x"580000",x"400000",x"2c2c2c",
x"484848",x"bc0000",x"640000",x"b4b4b4",x"b4b4b4",x"7c0000",x"b4b4b4",x"989898",x"989898",x"707070",x"484848",x"580058",x"500050",x"480048",x"480048",x"480048",x"500050",x"480048",x"500050",x"580058",x"6c0070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"646464",x"6c0070",x"9c009c",x"6c0070",x"6c0070",x"9c009c",x"6c0070",x"646464",x"500050",x"500050",x"580058",x"580058",x"580058",x"580058",x"580058",x"840084",x"580058",x"580058",x"500050",x"480048",x"480048",x"480048",x"400040",x"400040",x"400040",x"484848",x"707070",x"989898",x"989898",x"b4b4b4",x"880000",x"b4b4b4",x"b4b4b4",x"580000",x"400000",x"2c2c2c",
x"484848",x"bc0000",x"b00000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"500050",x"580058",x"484848",x"646464",x"707070",x"707070",x"646464",x"646464",x"545454",x"484848",x"404040",x"303030",x"480048",x"500050",x"580058",x"840084",x"580058",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"9c009c",x"6c0070",x"6c0070",x"6c0070",x"6c0070",x"9c009c",x"7c7c7c",x"500050",x"580058",x"500050",x"580058",x"580058",x"840084",x"580058",x"580058",x"580058",x"545454",x"545454",x"484848",x"404040",x"383838",x"404040",x"484848",x"545454",x"646464",x"484848",x"600064",x"6c0070",x"c0c0c0",x"980000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"545454",x"bc0000",x"700000",x"a8a8a8",x"a8a8a8",x"700000",x"a8a8a8",x"500050",x"500050",x"580058",x"580058",x"580058",x"580058",x"500050",x"480048",x"500050",x"480048",x"500050",x"480048",x"500050",x"480048",x"500050",x"580058",x"840084",x"6c0070",x"500050",x"500050",x"500050",x"545454",x"6c0070",x"6c0070",x"6c0070",x"6c0070",x"6c0070",x"6c0070",x"545454",x"500050",x"500050",x"580058",x"6c0070",x"840084",x"580058",x"580058",x"580058",x"580058",x"500050",x"480048",x"480048",x"480048",x"480048",x"400040",x"480048",x"480048",x"500050",x"580058",x"600064",x"6c0070",x"d0d0d0",x"980000",x"d0d0d0",x"d0d0d0",x"580000",x"400000",x"2c2c2c",
x"484848",x"c80000",x"a40000",x"a8a8a8",x"a8a8a8",x"640000",x"a8a8a8",x"500050",x"500050",x"500050",x"580058",x"580058",x"580058",x"500050",x"500050",x"480048",x"500050",x"480048",x"500050",x"480048",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"9c009c",x"6c0070",x"6c0070",x"6c0070",x"6c0070",x"9c009c",x"7c7c7c",x"500050",x"580058",x"500050",x"580058",x"500050",x"580058",x"580058",x"580058",x"500050",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"500050",x"580058",x"580058",x"600064",x"600064",x"c0c0c0",x"980000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"484848",x"a40000",x"980000",x"989898",x"989898",x"4c0000",x"989898",x"500050",x"500050",x"580058",x"500050",x"580058",x"500050",x"580058",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"6c0070",x"9c009c",x"484848",x"6c0070",x"9c009c",x"6c0070",x"545454",x"500050",x"500050",x"580058",x"500050",x"580058",x"580058",x"580058",x"500050",x"500050",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"500050",x"500050",x"600064",x"6c0070",x"600064",x"c0c0c0",x"880000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"484848",x"484848",x"383838",x"a8a8a8",x"a8a8a8",x"580000",x"a8a8a8",x"500050",x"500050",x"500050",x"580058",x"500050",x"580058",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"500050",x"500050",x"500050",x"500050",x"545454",x"500050",x"500050",x"500050",x"7c7c7c",x"545454",x"6c0070",x"484848",x"6c0070",x"6c0070",x"545454",x"7c7c7c",x"500050",x"580058",x"500050",x"545454",x"580058",x"500050",x"500050",x"500050",x"545454",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"480048",x"500050",x"500050",x"600064",x"600064",x"500050",x"b4b4b4",x"7c0000",x"b4b4b4",x"b4b4b4",x"202020",x"202020",x"2c2c2c",
x"545454",x"545454",x"545454",x"a8a8a8",x"a8a8a8",x"640000",x"a8a8a8",x"646464",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"484848",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"500050",x"500050",x"500050",x"500050",x"545454",x"7c7c7c",x"7c7c7c",x"545454",x"545454",x"7c7c7c",x"7c7c7c",x"545454",x"500050",x"500050",x"500050",x"580058",x"545454",x"500050",x"500050",x"480048",x"500050",x"480048",x"707070",x"484848",x"480048",x"480048",x"480048",x"500050",x"500050",x"580058",x"600064",x"580058",x"646464",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"2c2c2c",x"2c2c2c",
x"bc0000",x"bc0000",x"bc0000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"989898",x"646464",x"500050",x"500050",x"500050",x"500050",x"484848",x"707070",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"7c7c7c",x"7c7c7c",x"545454",x"500050",x"500050",x"500050",x"500050",x"580058",x"500050",x"500050",x"707070",x"500050",x"500050",x"480048",x"480048",x"480048",x"500050",x"707070",x"707070",x"484848",x"500050",x"500050",x"580058",x"580058",x"646464",x"989898",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"bc0000",
x"a40000",x"b00000",x"a40000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"989898",x"989898",x"989898",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"480048",x"500050",x"480048",x"480048",x"480048",x"480048",x"500050",x"707070",x"989898",x"989898",x"989898",x"989898",x"b4b4b4",x"a8a8a8",x"a8a8a8",x"640000",x"a8a8a8",x"a8a8a8",x"580000",x"580000",x"a40000",
x"a40000",x"7c0000",x"880000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"989898",x"989898",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"480048",x"500050",x"480048",x"500050",x"480048",x"500050",x"580058",x"580058",x"580058",x"707070",x"989898",x"989898",x"989898",x"989898",x"580000",x"989898",x"989898",x"580000",x"580000",x"700000",
x"880000",x"7c0000",x"a40000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"707070",x"480048",x"500050",x"480048",x"500050",x"580058",x"580058",x"580058",x"580058",x"580058",x"500050",x"500050",x"8c8c8c",x"8c8c8c",x"4c0000",x"8c8c8c",x"8c8c8c",x"580000",x"580000",x"700000",
x"a40000",x"880000",x"7c0000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"646464",x"989898",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"989898",x"646464",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"580058",x"580058",x"580058",x"580058",x"500050",x"500050",x"989898",x"989898",x"580000",x"989898",x"989898",x"580000",x"580000",x"880000",
x"a40000",x"880000",x"7c0000",x"b4b4b4",x"b4b4b4",x"7c0000",x"b4b4b4",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"580058",x"580058",x"580058",x"580058",x"580058",x"500050",x"707070",x"989898",x"989898",x"640000",x"989898",x"989898",x"580000",x"580000",x"700000",
x"700000",x"700000",x"880000",x"b4b4b4",x"b4b4b4",x"7c0000",x"b4b4b4",x"b4b4b4",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"580058",x"500050",x"580058",x"500050",x"500050",x"989898",x"a8a8a8",x"a8a8a8",x"640000",x"a8a8a8",x"a8a8a8",x"580000",x"580000",x"700000",
x"400000",x"400000",x"4c0000",x"b4b4b4",x"b4b4b4",x"880000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"580058",x"500050",x"707070",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"640000",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"400000",
x"2c2c2c",x"2c2c2c",x"2c2c2c",x"c0c0c0",x"c0c0c0",x"880000",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"707070",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"202020",x"2c2c2c",
x"545454",x"484848",x"545454",x"d0d0d0",x"d0d0d0",x"a40000",x"d0d0d0",x"d0d0d0",x"d0d0d0",x"b4b4b4",x"b4b4b4",x"989898",x"989898",x"989898",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"b4b4b4",x"9c009c",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"9c009c",x"b4b4b4",x"989898",x"500050",x"500050",x"500050",x"500050",x"500050",x"989898",x"989898",x"989898",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"2c2c2c",x"2c2c2c",
x"383838",x"ec0000",x"d40000",x"c0c0c0",x"c0c0c0",x"980000",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"989898",x"500050",x"500050",x"500050",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"707070",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"707070",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"500050",x"500050",x"500050",x"989898",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"880000",x"c0c0c0",x"c0c0c0",x"580000",x"580000",x"2c2c2c",
x"545454",x"d40000",x"a40000",x"b4b4b4",x"b4b4b4",x"980000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"b45400",x"b45400",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"b45400",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b45400",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"b45400",x"b45400",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"880000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"484848",x"d40000",x"a40000",x"b4b4b4",x"b4b4b4",x"880000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"744c28",x"744c28",x"500050",x"500050",x"707070",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"707070",x"500050",x"500050",x"744c28",x"744c28",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"d0d0d0",x"d0d0d0",x"d0d0d0",x"980000",x"d0d0d0",x"d0d0d0",x"580000",x"400000",x"2c2c2c",
x"484848",x"d40000",x"880000",x"b4b4b4",x"b4b4b4",x"880000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"646464",x"744c28",x"b45400",x"b45400",x"b45400",x"b45400",x"744c28",x"744c28",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"744c28",x"744c28",x"b45400",x"b45400",x"b45400",x"b45400",x"744c28",x"646464",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"980000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"383838",x"d40000",x"a40000",x"b4b4b4",x"b4b4b4",x"7c0000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"b45400",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"c0c0c0",x"c0c0c0",x"880000",x"c0c0c0",x"c0c0c0",x"580000",x"400000",x"2c2c2c",
x"545454",x"d40000",x"a40000",x"a8a8a8",x"a8a8a8",x"700000",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b45400",x"744c28",x"744c28",x"8c8c8c",x"b45400",x"b45400",x"744c28",x"b4b4b4",x"8c8c8c",x"744c28",x"b45400",x"b4b4b4",x"7c7c7c",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"b4b4b4",x"b45400",x"744c28",x"8c8c8c",x"b4b4b4",x"744c28",x"b45400",x"b45400",x"8c8c8c",x"744c28",x"744c28",x"b45400",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"400000",x"2c2c2c",
x"383838",x"c80000",x"a40000",x"a8a8a8",x"a8a8a8",x"700000",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"b4b4b4",x"744c28",x"7c7c7c",x"8c8c8c",x"b4b4b4",x"b45400",x"744c28",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"744c28",x"b45400",x"b4b4b4",x"8c8c8c",x"7c7c7c",x"744c28",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"580000",x"400000",x"2c2c2c",
x"545454",x"a40000",x"640000",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b45400",x"744c28",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"744c28",x"b45400",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"700000",x"b4b4b4",x"b4b4b4",x"400000",x"400000",x"2c2c2c",
x"383838",x"484848",x"2c2c2c",x"b4b4b4",x"b4b4b4",x"700000",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"b45400",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b45400",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"202020",x"2c2c2c",
x"545454",x"383838",x"545454",x"b4b4b4",x"b4b4b4",x"700000",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"500050",x"500050",x"500050",x"500050",x"500050",x"646464",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"646464",x"500050",x"500050",x"500050",x"500050",x"500050",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"700000",x"b4b4b4",x"b4b4b4",x"202020",x"2c2c2c",x"2c2c2c",
x"d40000",x"d40000",x"d40000",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"500050",x"500050",x"646464",x"b4b4b4",x"7c7c7c",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"7c7c7c",x"b4b4b4",x"646464",x"500050",x"500050",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"580000",x"580000",x"bc0000",
x"7c0000",x"a40000",x"580000",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"8c8c8c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"7c7c7c",x"580000",x"580000",x"700000",
x"a40000",x"7c0000",x"7c0000",x"580000",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"500050",x"500050",x"500050",x"500050",x"500050",x"500050",x"646464",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"700000",x"8c8c8c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"580000",x"580000",x"580000",x"4c0000",
x"a40000",x"7c0000",x"580000",x"580000",x"580000",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"500050",x"500050",x"500050",x"500050",x"646464",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"580000",x"580000",x"580000",x"700000",x"880000",
x"7c0000",x"980000",x"580000",x"580000",x"580000",x"580000",x"580000",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"500050",x"500050",x"646464",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"580000",x"580000",x"580000",x"580000",x"580000",x"640000",x"700000",x"a40000",
x"640000",x"a40000",x"7c0000",x"a40000",x"640000",x"580000",x"640000",x"580000",x"580000",x"580000",x"580000",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"646464",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"580000",x"580000",x"580000",x"580000",x"580000",x"580000",x"700000",x"580000",x"a40000",x"700000",x"a40000",
x"640000",x"a40000",x"7c0000",x"7c0000",x"640000",x"980000",x"980000",x"640000",x"580000",x"580000",x"580000",x"580000",x"580000",x"580000",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"580000",x"580000",x"580000",x"580000",x"580000",x"580000",x"580000",x"700000",x"a40000",x"700000",x"580000",x"640000",x"a40000",x"4c0000",
x"7c0000",x"980000",x"580000",x"a40000",x"640000",x"640000",x"880000",x"640000",x"7c0000",x"7c0000",x"a40000",x"580000",x"580000",x"580000",x"580000",x"580000",x"580000",x"400000",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"400000",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"580000",x"580000",x"580000",x"580000",x"a40000",x"580000",x"a40000",x"700000",x"a40000",x"700000",x"a40000",x"640000",x"a40000",x"700000",
x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"400000",x"400000",x"202020",x"202020",x"2c2c2c",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"989898",x"7c7c7c",x"700000",x"700000",x"700000",x"700000",x"7c7c7c",x"989898",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"4c0000",x"4c0000",x"4c0000",x"400000",x"400000",x"202020",x"2c2c2c",x"2c2c2c",x"580000",x"400000",x"400000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",x"4c0000",
x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",
x"383838",x"545454",x"383838",x"545454",x"383838",x"383838",x"383838",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"545454",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"7c7c7c",x"545454",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"383838",x"484848",x"484848",x"545454",x"484848",x"484848",x"484848",x"484848",x"404040",x"383838",x"404040",x"484848",x"484848",x"484848",
x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"383838",x"383838",x"383838",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",


--10 colorstone



x"7c7c7c",x"7c7c7c",x"7c7c7c",x"483818",x"543c1c",x"5c4020",x"5c4020",x"744c28",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"483818",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"483818",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"707070",x"707070",x"707070",x"707070",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"484848",x"646464",x"707070",x"545454",x"646464",x"545454",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"545454",x"5c5c5c",x"5c5c5c",x"646464",x"707070",x"7c7c7c",
x"7c7c7c",x"707070",x"707070",x"545454",x"483818",x"543c1c",x"5c4020",x"744c28",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"483818",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"483818",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"707070",x"7c7c7c",x"707070",x"7c7c7c",x"7c7c7c",x"484848",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"484848",x"646464",x"707070",x"545454",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"545454",x"545454",x"5c5c5c",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"707070",
x"707070",x"707070",x"707070",x"646464",x"545454",x"483818",x"543c1c",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"483818",x"5c4020",x"543c1c",x"543c1c",x"483818",x"484848",x"545454",x"646464",x"646464",x"484848",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"484848",x"646464",x"646464",x"484848",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"484848",x"646464",x"707070",x"545454",x"646464",x"545454",x"4c4c4c",x"545454",x"5c5c5c",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",
x"545454",x"707070",x"7c7c7c",x"707070",x"646464",x"545454",x"483818",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"403018",x"483818",x"543c1c",x"483818",x"483818",x"545454",x"646464",x"7c7c7c",x"484848",x"5c4020",x"5c4020",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"646464",x"646464",x"484848",x"484848",x"484848",x"646464",x"707070",x"545454",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"5c5c5c",x"545454",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"545454",x"707070",x"707070",x"7c7c7c",x"646464",x"483818",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"403018",x"483818",x"483818",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"484848",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"484848",x"7c7c7c",x"646464",x"646464",x"646464",x"707070",x"545454",x"646464",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"5c5c5c",
x"4c4c4c",x"4c4c4c",x"545454",x"707070",x"707070",x"707070",x"483818",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"403018",x"483818",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"5c4020",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"403018",x"382c14",x"646464",x"8c8c8c",x"a8a8a8",x"707070",x"545454",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"545454",x"707070",x"7c7c7c",x"545454",x"483818",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"403018",x"484848",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"484848",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"483818",x"382c14",x"382c14",x"646464",x"a8a8a8",x"7c7c7c",x"545454",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"545454",x"707070",x"7c7c7c",x"545454",x"483818",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"403018",x"483818",x"545454",x"646464",x"646464",x"7c7c7c",x"646464",x"5c4020",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"483818",x"382c14",x"382c14",x"646464",x"989898",x"7c7c7c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"545454",x"7c7c7c",x"646464",x"545454",x"483818",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"403018",x"403018",x"545454",x"646464",x"646464",x"7c7c7c",x"7c7c7c",x"484848",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"483818",x"403018",x"382c14",x"483818",x"382c14",x"382c14",x"646464",x"989898",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"483818",x"543c1c",x"543c1c",x"543c1c",x"543c1c",x"403018",x"403018",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"646464",x"5c4020",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"483818",x"403018",x"382c14",x"403018",x"382c14",x"382c14",x"646464",x"8c8c8c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"7c7c7c",x"707070",x"7c7c7c",x"646464",x"545454",x"403018",x"403018",x"403018",x"403018",x"484848",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"484848",x"5c4020",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"403018",x"382c14",x"404040",x"646464",x"8c8c8c",x"646464",x"5c5c5c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"707070",x"707070",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"5c4020",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"382c14",x"4c4c4c",x"707070",x"7c7c7c",x"646464",x"5c5c5c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"383838",x"707070",x"707070",x"646464",x"545454",x"545454",x"545454",x"646464",x"707070",x"989898",x"989898",x"8c8c8c",x"707070",x"646464",x"5c4020",x"543c1c",x"543c1c",x"483818",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"382c14",x"545454",x"707070",x"8c8c8c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"4c4c4c",x"484848",x"484848",x"484848",x"484848",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"383838",x"646464",x"7c7c7c",x"646464",x"545454",x"545454",x"545454",x"545454",x"484848",x"646464",x"989898",x"8c8c8c",x"8c8c8c",x"646464",x"5c4020",x"483818",x"543c1c",x"543c1c",x"483818",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"382c14",x"646464",x"707070",x"7c7c7c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"484848",x"484848",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"4c4c4c",x"484848",x"383838",x"646464",x"7c7c7c",x"707070",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"707070",x"8c8c8c",x"7c7c7c",x"5c4020",x"543c1c",x"483818",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"404040",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"484848",x"484848",x"4c4c4c",x"4c4c4c",
x"4c4c4c",x"484848",x"383838",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"646464",x"545454",x"5c4020",x"483818",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"4c4c4c",x"707070",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"484848",x"484848",x"484848",x"4c4c4c",x"484848",
x"484848",x"383838",x"646464",x"7c7c7c",x"7c7c7c",x"707070",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"404040",x"4c4c4c",x"545454",x"484848",x"646464",x"5c4020",x"483818",x"5c4020",x"483818",x"483818",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"483818",x"483818",x"403018",x"382c14",x"382c14",x"545454",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"383838",
x"383838",x"646464",x"646464",x"484848",x"484848",x"646464",x"707070",x"545454",x"545454",x"545454",x"545454",x"4c4c4c",x"404040",x"545454",x"545454",x"646464",x"646464",x"5c4020",x"483818",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"483818",x"483818",x"403018",x"382c14",x"382c14",x"646464",x"6c4824",x"5c4020",x"646464",x"545454",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"383838",x"404040",
x"646464",x"646464",x"484848",x"543c1c",x"543c1c",x"484848",x"646464",x"646464",x"545454",x"545454",x"545454",x"404040",x"404040",x"545454",x"545454",x"545454",x"707070",x"5c4020",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"403018",x"483818",x"403018",x"382c14",x"403018",x"5c5c5c",x"6c4824",x"5c4020",x"5c4020",x"545454",x"646464",x"404040",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"404040",x"383838",x"404040",x"404040",
x"646464",x"484848",x"543c1c",x"5c4020",x"483818",x"543c1c",x"484848",x"7c7c7c",x"484848",x"545454",x"404040",x"404040",x"404040",x"545454",x"545454",x"545454",x"646464",x"646464",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"403018",x"382c14",x"382c14",x"403018",x"646464",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"646464",x"404040",x"484848",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"404040",x"383838",x"343434",x"343434",x"383838",x"404040",x"646464",
x"484848",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"403018",x"646464",x"707070",x"484848",x"404040",x"545454",x"404040",x"545454",x"545454",x"545454",x"484848",x"7c7c7c",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"382c14",x"382c14",x"382c14",x"4c4c4c",x"646464",x"7c7c7c",x"483818",x"483818",x"483818",x"483818",x"483818",x"707070",x"707070",x"646464",x"404040",x"404040",x"404040",x"484848",x"484848",x"484848",x"484848",x"484848",x"404040",x"404040",x"383838",x"343434",x"383838",x"404040",x"383838",x"545454",x"646464",x"646464",
x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"403018",x"484848",x"7c7c7c",x"646464",x"484848",x"545454",x"404040",x"545454",x"545454",x"545454",x"484848",x"707070",x"646464",x"403018",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"382c14",x"382c14",x"4c4c4c",x"646464",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"646464",x"646464",x"646464",x"646464",x"8c8c8c",x"8c8c8c",x"646464",x"646464",x"404040",x"383838",x"343434",x"343434",x"343434",x"343434",x"343434",x"343434",x"343434",x"383838",x"404040",x"404040",x"383838",x"545454",x"646464",x"7c7c7c",x"484848",
x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"646464",x"707070",x"484848",x"545454",x"404040",x"545454",x"545454",x"545454",x"383838",x"646464",x"7c7c7c",x"484848",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"382c14",x"404040",x"5c5c5c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"7c7c7c",x"8c8c8c",x"989898",x"989898",x"707070",x"646464",x"545454",x"383838",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"383838",x"545454",x"646464",x"7c7c7c",x"484848",x"543c1c",
x"483818",x"483818",x"483818",x"543c1c",x"483818",x"483818",x"403018",x"483818",x"646464",x"7c7c7c",x"646464",x"484848",x"404040",x"545454",x"545454",x"4c4c4c",x"383838",x"646464",x"7c7c7c",x"646464",x"403018",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"382c14",x"404040",x"545454",x"646464",x"646464",x"545454",x"484848",x"404040",x"383838",x"404040",x"404040",x"404040",x"404040",x"545454",x"7c7c7c",x"989898",x"989898",x"8c8c8c",x"7c7c7c",x"646464",x"545454",x"383838",x"404040",x"404040",x"404040",x"404040",x"404040",x"383838",x"383838",x"545454",x"646464",x"7c7c7c",x"484848",x"543c1c",x"5c4020",
x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"484848",x"7c7c7c",x"7c7c7c",x"646464",x"404040",x"545454",x"4c4c4c",x"484848",x"383838",x"646464",x"7c7c7c",x"7c7c7c",x"484848",x"382c14",x"403018",x"483818",x"483818",x"483818",x"403018",x"382c14",x"382c14",x"545454",x"646464",x"7c7c7c",x"646464",x"545454",x"484848",x"404040",x"404040",x"383838",x"383838",x"404040",x"404040",x"404040",x"404040",x"545454",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"707070",x"7c7c7c",x"646464",x"545454",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"545454",x"646464",x"7c7c7c",x"646464",x"543c1c",x"5c4020",x"483818",
x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"646464",x"7c7c7c",x"707070",x"383838",x"484848",x"484848",x"484848",x"383838",x"707070",x"707070",x"7c7c7c",x"646464",x"382c14",x"382c14",x"382c14",x"382c14",x"382c14",x"382c14",x"382c14",x"404040",x"646464",x"7c7c7c",x"646464",x"545454",x"484848",x"404040",x"404040",x"404040",x"383838",x"404040",x"383838",x"404040",x"404040",x"383838",x"404040",x"707070",x"7c7c7c",x"707070",x"545454",x"545454",x"7c7c7c",x"646464",x"545454",x"383838",x"383838",x"383838",x"383838",x"545454",x"646464",x"7c7c7c",x"646464",x"484848",x"5c4020",x"483818",x"483818",
x"483818",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"382c14",x"483818",x"403018",x"545454",x"707070",x"7c7c7c",x"646464",x"383838",x"383838",x"383838",x"707070",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"484848",x"382c14",x"382c14",x"382c14",x"382c14",x"404040",x"4c4c4c",x"5c5c5c",x"7c7c7c",x"545454",x"545454",x"484848",x"404040",x"484848",x"484848",x"404040",x"383838",x"404040",x"383838",x"404040",x"404040",x"383838",x"484848",x"646464",x"707070",x"646464",x"484848",x"484848",x"545454",x"7c7c7c",x"646464",x"545454",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"483818",
x"483818",x"543c1c",x"543c1c",x"483818",x"483818",x"483818",x"382c14",x"483818",x"403018",x"484848",x"7c7c7c",x"8c8c8c",x"707070",x"646464",x"646464",x"707070",x"7c7c7c",x"545454",x"6c4824",x"6c4824",x"545454",x"646464",x"484848",x"484848",x"4c4c4c",x"5c5c5c",x"5c5c5c",x"7c7c7c",x"7c7c7c",x"545454",x"545454",x"484848",x"404040",x"404040",x"484848",x"484848",x"404040",x"383838",x"404040",x"404040",x"383838",x"404040",x"343434",x"545454",x"646464",x"707070",x"545454",x"484848",x"484848",x"484848",x"545454",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"707070",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"483818",x"543c1c",x"483818",x"483818",x"382c14",x"483818",x"403018",x"484848",x"7c7c7c",x"707070",x"8c8c8c",x"707070",x"707070",x"646464",x"6c4824",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"646464",x"646464",x"646464",x"707070",x"7c7c7c",x"707070",x"545454",x"545454",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"343434",x"404040",x"404040",x"383838",x"383838",x"303030",x"545454",x"646464",x"646464",x"484848",x"484848",x"484848",x"484848",x"484848",x"646464",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"707070",x"646464",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"483818",x"403018",x"484848",x"7c7c7c",x"707070",x"707070",x"707070",x"707070",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"7c7c7c",x"7c7c7c",x"707070",x"707070",x"545454",x"545454",x"484848",x"404040",x"404040",x"404040",x"484848",x"404040",x"404040",x"404040",x"343434",x"404040",x"404040",x"383838",x"383838",x"484848",x"646464",x"707070",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"545454",x"646464",x"707070",x"707070",x"646464",x"5c5c5c",x"545454",x"543c1c",x"483818",x"483818",x"543c1c",x"543c1c",x"543c1c",
x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"483818",x"403018",x"545454",x"707070",x"8c8c8c",x"707070",x"707070",x"707070",x"646464",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"7c7c7c",x"707070",x"7c7c7c",x"545454",x"545454",x"545454",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"343434",x"404040",x"404040",x"383838",x"343434",x"545454",x"707070",x"7c7c7c",x"7c7c7c",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"7c7c7c",x"707070",x"5c5c5c",x"545454",x"5c5c5c",x"543c1c",x"483818",x"483818",x"543c1c",x"543c1c",x"543c1c",
x"483818",x"483818",x"483818",x"483818",x"483818",x"382c14",x"403018",x"403018",x"403018",x"545454",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"483818",x"7c7c7c",x"7c7c7c",x"545454",x"545454",x"484848",x"545454",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"343434",x"404040",x"404040",x"383838",x"303030",x"646464",x"545454",x"744c28",x"744c28",x"744c28",x"744c28",x"744c28",x"744c28",x"744c28",x"744c28",x"744c28",x"483818",x"5c4020",x"744c28",x"5c5c5c",x"646464",x"543c1c",x"483818",x"483818",x"543c1c",x"543c1c",x"543c1c",
x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"483818",x"403018",x"484848",x"646464",x"7c7c7c",x"646464",x"545454",x"5c5c5c",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"543c1c",x"543c1c",x"483818",x"483818",x"646464",x"7c7c7c",x"545454",x"545454",x"484848",x"484848",x"545454",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"404040",x"404040",x"343434",x"545454",x"707070",x"6c4824",x"6c4824",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"5c4020",x"5c4020",x"5c4020",x"7c7c7c",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"483818",x"483818",x"403018",x"382c14",x"403018",x"484848",x"646464",x"646464",x"646464",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"545454",x"7c7c7c",x"646464",x"545454",x"484848",x"404040",x"484848",x"545454",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"383838",x"303030",x"404040",x"383838",x"303030",x"545454",x"646464",x"6c4824",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"5c4020",x"5c4020",x"543c1c",x"646464",x"543c1c",x"483818",x"483818",x"543c1c",x"483818",x"483818",
x"483818",x"483818",x"483818",x"483818",x"382c14",x"403018",x"484848",x"646464",x"646464",x"7c7c7c",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"545454",x"484848",x"404040",x"404040",x"484848",x"545454",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"383838",x"303030",x"404040",x"383838",x"303030",x"646464",x"545454",x"80502c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"5c4020",x"5c4020",x"543c1c",x"646464",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"483818",x"403018",x"382c14",x"484848",x"646464",x"646464",x"707070",x"646464",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"545454",x"404040",x"404040",x"404040",x"484848",x"545454",x"4c4c4c",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"343434",x"303030",x"404040",x"303030",x"646464",x"707070",x"484848",x"80502c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"5c4020",x"5c4020",x"543c1c",x"646464",x"403018",x"483818",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"483818",x"382c14",x"484848",x"646464",x"646464",x"7c7c7c",x"7c7c7c",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"8c8c8c",x"989898",x"989898",x"545454",x"404040",x"404040",x"404040",x"484848",x"545454",x"4c4c4c",x"404040",x"404040",x"404040",x"404040",x"404040",x"404040",x"343434",x"303030",x"383838",x"484848",x"707070",x"707070",x"6c4824",x"80502c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"5c4020",x"5c4020",x"543c1c",x"646464",x"484848",x"403018",x"483818",x"483818",x"483818",x"483818",
x"483818",x"483818",x"403018",x"484848",x"646464",x"646464",x"707070",x"7c7c7c",x"646464",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"989898",x"989898",x"646464",x"404040",x"404040",x"404040",x"484848",x"545454",x"4c4c4c",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"303030",x"343434",x"545454",x"7c7c7c",x"646464",x"6c4824",x"80502c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"543c1c",x"646464",x"646464",x"484848",x"403018",x"483818",x"483818",x"483818",
x"483818",x"403018",x"484848",x"646464",x"646464",x"707070",x"7c7c7c",x"646464",x"545454",x"5c5c5c",x"545454",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"545454",x"646464",x"8c8c8c",x"707070",x"383838",x"404040",x"404040",x"484848",x"545454",x"4c4c4c",x"484848",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"303030",x"303030",x"646464",x"7c7c7c",x"545454",x"6c4824",x"80502c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"543c1c",x"646464",x"7c7c7c",x"646464",x"484848",x"403018",x"483818",x"483818",
x"403018",x"484848",x"646464",x"646464",x"7c7c7c",x"7c7c7c",x"707070",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"545454",x"8c8c8c",x"8c8c8c",x"545454",x"383838",x"383838",x"484848",x"545454",x"484848",x"4c4c4c",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"303030",x"484848",x"707070",x"707070",x"6c4824",x"5c4020",x"80502c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"484848",x"403018",x"403018",
x"484848",x"646464",x"646464",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"404040",x"545454",x"545454",x"646464",x"707070",x"707070",x"303030",x"383838",x"383838",x"545454",x"404040",x"4c4c4c",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"303030",x"545454",x"7c7c7c",x"646464",x"6c4824",x"5c4020",x"80502c",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"646464",x"484848",x"484848",
x"646464",x"646464",x"989898",x"989898",x"8c8c8c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"404040",x"484848",x"545454",x"545454",x"646464",x"646464",x"484848",x"303030",x"343434",x"303030",x"404040",x"4c4c4c",x"404040",x"404040",x"404040",x"404040",x"404040",x"303030",x"303030",x"545454",x"7c7c7c",x"545454",x"6c4824",x"5c4020",x"80502c",x"744c28",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"383838",x"545454",x"646464",x"646464",
x"646464",x"7c7c7c",x"989898",x"989898",x"707070",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"484848",x"404040",x"545454",x"545454",x"545454",x"646464",x"545454",x"484848",x"303030",x"303030",x"383838",x"484848",x"484848",x"404040",x"404040",x"404040",x"383838",x"303030",x"484848",x"646464",x"707070",x"6c4824",x"5c4020",x"5c4020",x"744c28",x"80502c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"545454",
x"2c2c2c",x"484848",x"8c8c8c",x"8c8c8c",x"646464",x"545454",x"545454",x"545454",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"404040",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"646464",x"545454",x"343434",x"343434",x"484848",x"404040",x"404040",x"404040",x"383838",x"303030",x"545454",x"707070",x"7c7c7c",x"6c4824",x"5c4020",x"5c4020",x"6c4824",x"80502c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"2c2c2c",
x"2c2c2c",x"202020",x"484848",x"7c7c7c",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"484848",x"404040",x"484848",x"545454",x"545454",x"545454",x"484848",x"646464",x"646464",x"545454",x"303030",x"343434",x"343434",x"383838",x"404040",x"404040",x"383838",x"303030",x"646464",x"7c7c7c",x"7c7c7c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"744c28",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"2c2c2c",
x"2c2c2c",x"202020",x"484848",x"707070",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"404040",x"484848",x"545454",x"545454",x"484848",x"383838",x"646464",x"8c8c8c",x"8c8c8c",x"545454",x"303030",x"343434",x"343434",x"404040",x"404040",x"343434",x"484848",x"707070",x"707070",x"707070",x"646464",x"543c1c",x"5c4020",x"5c4020",x"6c4824",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"2c2c2c",
x"202020",x"484848",x"646464",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"484848",x"404040",x"484848",x"545454",x"484848",x"383838",x"484848",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"545454",x"303030",x"343434",x"383838",x"383838",x"303030",x"545454",x"7c7c7c",x"707070",x"707070",x"7c7c7c",x"646464",x"543c1c",x"5c4020",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"543c1c",x"483818",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"2c2c2c",x"2c2c2c",
x"484848",x"646464",x"646464",x"646464",x"484848",x"545454",x"545454",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"484848",x"343434",x"484848",x"484848",x"383838",x"484848",x"545454",x"7c7c7c",x"484848",x"483818",x"484848",x"7c7c7c",x"545454",x"303030",x"303030",x"303030",x"303030",x"707070",x"7c7c7c",x"646464",x"383838",x"383838",x"646464",x"646464",x"543c1c",x"543c1c",x"5c4020",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"543c1c",x"483818",x"484848",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"2c2c2c",x"2c2c2c",
x"646464",x"707070",x"707070",x"707070",x"646464",x"484848",x"545454",x"5c5c5c",x"5c5c5c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"484848",x"343434",x"404040",x"383838",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"403018",x"484848",x"7c7c7c",x"646464",x"545454",x"545454",x"646464",x"7c7c7c",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"707070",x"646464",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"484848",x"646464",x"646464",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",
x"7c7c7c",x"7c7c7c",x"707070",x"707070",x"7c7c7c",x"646464",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"545454",x"404040",x"343434",x"383838",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"403018",x"483818",x"403018",x"484848",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"707070",x"646464",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"484848",x"646464",x"707070",x"7c7c7c",x"7c7c7c",x"484848",x"484848",x"484848",x"484848",x"484848",
x"7c7c7c",x"707070",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"646464",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"545454",x"404040",x"343434",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"484848",x"7c7c7c",x"7c7c7c",x"484848",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"707070",x"707070",x"545454",x"543c1c",x"543c1c",x"543c1c",x"483818",x"483818",x"484848",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"646464",x"7c7c7c",x"7c7c7c",
x"7c7c7c",x"545454",x"6c4824",x"6c4824",x"545454",x"8c8c8c",x"8c8c8c",x"646464",x"484848",x"383838",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"343434",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"403018",x"7c7c7c",x"646464",x"383838",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"707070",x"545454",x"543c1c",x"483818",x"484848",x"484848",x"646464",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"646464",x"7c7c7c",
x"6c4824",x"6c4824",x"5c4020",x"5c4020",x"6c4824",x"6c4824",x"545454",x"7c7c7c",x"646464",x"484848",x"383838",x"484848",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"383838",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"403018",x"7c7c7c",x"383838",x"2c2c2c",x"2c2c2c",x"282828",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"707070",x"545454",x"484848",x"484848",x"646464",x"7c7c7c",x"545454",x"545454",x"545454",x"4c4c4c",x"545454",x"545454",x"545454",x"484848",x"646464",x"7c7c7c",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"6c4824",x"6c4824",x"545454",x"646464",x"484848",x"383838",x"484848",x"545454",x"484848",x"484848",x"383838",x"383838",x"484848",x"646464",x"484848",x"484848",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"483818",x"403018",x"403018",x"484848",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"707070",x"646464",x"646464",x"8c8c8c",x"646464",x"4c4c4c",x"4c4c4c",x"545454",x"545454",x"545454",x"545454",x"4c4c4c",x"484848",x"646464",x"7c7c7c",
x"5c4020",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"6c4824",x"483818",x"646464",x"484848",x"383838",x"484848",x"484848",x"383838",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"403018",x"484848",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"2c2c2c",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"707070",x"8c8c8c",x"8c8c8c",x"545454",x"4c4c4c",x"4c4c4c",x"545454",x"545454",x"545454",x"545454",x"4c4c4c",x"484848",x"646464",x"6c4824",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"483818",x"5c4020",x"5c4020",x"484848",x"383838",x"383838",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"403018",x"403018",x"545454",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"8c8c8c",x"646464",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"4c4c4c",x"484848",x"484848",x"646464",x"6c4824",
x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"483818",x"5c4020",x"5c4020",x"543c1c",x"484848",x"484848",x"545454",x"646464",x"484848",x"543c1c",x"543c1c",x"5c4020",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"403018",x"484848",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"545454",x"6c4824",x"5c4020",
x"5c4020",x"5c4020",x"543c1c",x"543c1c",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"5c4020",x"483818",x"543c1c",x"483818",x"483818",x"545454",x"545454",x"646464",x"484848",x"543c1c",x"483818",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"483818",x"403018",x"484848",x"646464",x"484848",x"383838",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"282828",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"202020",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"7c7c7c",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"4c4c4c",x"484848",x"646464",x"6c4824",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"543c1c",x"403018",x"483818",x"483818",x"545454",x"646464",x"646464",x"484848",x"543c1c",x"483818",x"483818",x"543c1c",x"5c4020",x"483818",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"403018",x"545454",x"646464",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"282828",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"646464",x"545454",x"545454",x"545454",x"4c4c4c",x"484848",x"484848",x"545454",x"6c4824",x"5c4020",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"483818",x"403018",x"483818",x"545454",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"484848",x"483818",x"483818",x"483818",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"403018",x"484848",x"646464",x"383838",x"2c2c2c",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"202020",x"282828",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"646464",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"484848",x"4c4c4c",x"484848",x"545454",x"6c4824",x"5c4020",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"403018",x"403018",x"545454",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"545454",x"483818",x"483818",x"483818",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"484848",x"646464",x"484848",x"383838",x"2c2c2c",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"202020",x"202020",x"282828",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"646464",x"4c4c4c",x"484848",x"545454",x"545454",x"484848",x"6c4824",x"5c4020",x"5c4020",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"483818",x"403018",x"403018",x"545454",x"7c7c7c",x"545454",x"404040",x"545454",x"7c7c7c",x"646464",x"484848",x"483818",x"483818",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"545454",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"1c1c1c",x"282828",x"282828",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"545454",x"646464",x"545454",x"545454",x"4c4c4c",x"646464",x"6c4824",x"5c4020",x"5c4020",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"483818",x"403018",x"545454",x"7c7c7c",x"545454",x"404040",x"404040",x"404040",x"545454",x"7c7c7c",x"545454",x"483818",x"483818",x"543c1c",x"5c4020",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"484848",x"646464",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"1c1c1c",x"202020",x"2c2c2c",x"202020",x"202020",x"282828",x"2c2c2c",x"2c2c2c",x"202020",x"545454",x"7c7c7c",x"4c4c4c",x"4c4c4c",x"646464",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",
x"5c4020",x"5c4020",x"5c4020",x"5c4020",x"543c1c",x"403018",x"403018",x"545454",x"7c7c7c",x"7c7c7c",x"404040",x"404040",x"404040",x"404040",x"404040",x"545454",x"646464",x"483818",x"483818",x"543c1c",x"483818",x"483818",x"483818",x"483818",x"483818",x"403018",x"484848",x"545454",x"646464",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"2c2c2c",x"2c2c2c",x"282828",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"282828",x"202020",x"1c1c1c",x"202020",x"2c2c2c",x"282828",x"202020",x"202020",x"282828",x"2c2c2c",x"202020",x"545454",x"7c7c7c",x"7c7c7c",x"646464",x"646464",x"6c4824",x"5c4020",x"5c4020",x"5c4020",x"5c4020",


--11 Mossy



x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",
x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"dcdcdc",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"b4ac00",x"b4ac00",x"b4ac00",x"dcdcdc",x"202020",x"383838",x"8c8c8c",x"a8a8a8",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"ccc400",x"ccc400",x"ccc400",x"707070",x"8c8c8c",x"8c8c8c",x"545454",x"202020",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",
x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"484848",x"dcdcdc",x"d0d0d0",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"989898",x"a8a8a8",x"ccc400",x"ccc400",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"ccc400",x"ccc400",x"8c8c8c",x"202020",x"383838",x"8c8c8c",x"c0c0c0",x"b4b4b4",x"8c8c8c",x"ccc400",x"7c7c7c",x"ccc400",x"9c9c00",x"9c9c00",x"9c9c00",x"706c00",x"545454",x"545454",x"383838",x"202020",x"383838",x"707070",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"707070",x"646464",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",
x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"202020",x"545454",x"484848",x"dcdcdc",x"d0d0d0",x"b4ac00",x"b4ac00",x"b4ac00",x"706c00",x"989898",x"ccc400",x"ccc400",x"9c9c00",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"848400",x"b4ac00",x"646464",x"202020",x"383838",x"a8a8a8",x"dcdcdc",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"ccc400",x"7c7c7c",x"706c00",x"848400",x"706c00",x"545454",x"7c7c7c",x"545454",x"383838",x"202020",x"383838",x"9c9c00",x"ccc400",x"e4d800",x"9c9c00",x"706c00",x"8c8c8c",x"b4b4b4",x"c0c0c0",x"ccc400",x"ccc400",x"ccc400",x"646464",x"646464",x"ccc400",x"ccc400",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",
x"d0d0d0",x"b4b4b4",x"b4ac00",x"b4b4b4",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"202020",x"545454",x"484848",x"dcdcdc",x"d0d0d0",x"9c9c00",x"9c9c00",x"848400",x"706c00",x"989898",x"ccc400",x"9c9c00",x"a8a8a8",x"a8a8a8",x"989898",x"8c8c8c",x"8c8c8c",x"9c9c00",x"545454",x"202020",x"383838",x"8c8c8c",x"c0c0c0",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"a8a8a8",x"646464",x"848400",x"706c00",x"545454",x"707070",x"545454",x"383838",x"202020",x"383838",x"9c9c00",x"e4d800",x"b4ac00",x"706c00",x"646464",x"7c7c7c",x"b4b4b4",x"dcdcdc",x"ccc400",x"e4d800",x"e4d800",x"484848",x"646464",x"ccc400",x"ccc400",x"848400",x"7c7c7c",x"d0d0d0",x"d0d0d0",
x"a8a8a8",x"a8a8a8",x"b4ac00",x"b4ac00",x"545454",x"707070",x"7c7c7c",x"707070",x"202020",x"545454",x"484848",x"dcdcdc",x"c0c0c0",x"9c9c00",x"848400",x"706c00",x"707070",x"7c7c7c",x"989898",x"a8a8a8",x"989898",x"9c9c00",x"8c8c8c",x"707070",x"8c8c8c",x"848400",x"545454",x"202020",x"383838",x"484848",x"a8a8a8",x"ccc400",x"9c9c00",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"585400",x"545454",x"707070",x"545454",x"545454",x"383838",x"202020",x"383838",x"9c9c00",x"e4d800",x"706c00",x"646464",x"8c8c8c",x"b4b4b4",x"e4d800",x"ccc400",x"7c7c7c",x"9c9c00",x"9c9c00",x"484848",x"646464",x"9c9c00",x"848400",x"706c00",x"484848",x"8c8c8c",x"989898",
x"b4b4b4",x"989898",x"706c00",x"545454",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"707070",x"202020",x"484848",x"484848",x"dcdcdc",x"d0d0d0",x"9c9c00",x"706c00",x"706c00",x"7c7c7c",x"a8a8a8",x"989898",x"989898",x"989898",x"9c9c00",x"8c8c8c",x"989898",x"707070",x"8c8c8c",x"545454",x"202020",x"383838",x"484848",x"7c7c7c",x"9c9c00",x"848400",x"b4ac00",x"8c8c8c",x"a8a8a8",x"a8a8a8",x"707070",x"646464",x"707070",x"383838",x"383838",x"383838",x"202020",x"383838",x"848400",x"9c9c00",x"706c00",x"646464",x"7c7c7c",x"ccc400",x"ccc400",x"ccc400",x"7c7c7c",x"706c00",x"9c9c00",x"484848",x"707070",x"646464",x"484848",x"484848",x"646464",x"b4ac00",x"7c7c7c",
x"b4b4b4",x"b4b4b4",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"707070",x"545454",x"202020",x"383838",x"484848",x"dcdcdc",x"d0d0d0",x"8c8c8c",x"7c7c7c",x"7c7c7c",x"989898",x"a8a8a8",x"989898",x"d0d0d0",x"7c7c7c",x"848400",x"989898",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"545454",x"202020",x"383838",x"484848",x"707070",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"707070",x"383838",x"383838",x"383838",x"2c2c2c",x"383838",x"848400",x"706c00",x"646464",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"ccc400",x"7c7c7c",x"7c7c7c",x"706c00",x"706c00",x"484848",x"707070",x"7c7c7c",x"8c8c8c",x"707070",x"7c7c7c",x"848400",x"646464",
x"989898",x"a8a8a8",x"a8a8a8",x"707070",x"707070",x"8c8c8c",x"484848",x"484848",x"202020",x"2c2c2c",x"484848",x"dcdcdc",x"c0c0c0",x"a8a8a8",x"989898",x"7c7c7c",x"989898",x"ccc400",x"989898",x"989898",x"8c8c8c",x"989898",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"545454",x"202020",x"202020",x"484848",x"545454",x"707070",x"707070",x"545454",x"545454",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"202020",x"383838",x"383838",x"7c7c7c",x"646464",x"8c8c8c",x"7c7c7c",x"a8a8a8",x"a8a8a8",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"7c7c7c",x"484848",x"707070",x"8c8c8c",x"989898",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"7c7c7c",x"646464",
x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"707070",x"545454",x"484848",x"484848",x"202020",x"2c2c2c",x"484848",x"dcdcdc",x"ececec",x"a8a8a8",x"7c7c7c",x"989898",x"7c7c7c",x"ccc400",x"b4ac00",x"707070",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"545454",x"2c2c2c",x"202020",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"202020",x"202020",x"383838",x"383838",x"383838",x"7c7c7c",x"b4b4b4",x"b4b4b4",x"8c8c8c",x"9c9c00",x"7c7c7c",x"989898",x"7c7c7c",x"7c7c7c",x"989898",x"646464",x"707070",x"989898",x"8c8c8c",x"989898",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",
x"707070",x"707070",x"707070",x"707070",x"545454",x"484848",x"383838",x"383838",x"202020",x"2c2c2c",x"484848",x"dcdcdc",x"dcdcdc",x"8c8c8c",x"7c7c7c",x"989898",x"989898",x"ccc400",x"9c9c00",x"707070",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"545454",x"2c2c2c",x"202020",x"383838",x"484848",x"383838",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"383838",x"383838",x"383838",x"383838",x"7c7c7c",x"b4b4b4",x"7c7c7c",x"9c9c00",x"484848",x"8c8c8c",x"a8a8a8",x"e4d800",x"7c7c7c",x"8c8c8c",x"707070",x"8c8c8c",x"707070",x"989898",x"646464",x"707070",x"8c8c8c",x"646464",x"646464",
x"545454",x"545454",x"484848",x"484848",x"484848",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"484848",x"a8a8a8",x"dcdcdc",x"a8a8a8",x"989898",x"7c7c7c",x"ccc400",x"b4ac00",x"9c9c00",x"707070",x"989898",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"707070",x"646464",x"383838",x"202020",x"383838",x"484848",x"484848",x"484848",x"484848",x"707070",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"dcdcdc",x"dcdcdc",x"706c00",x"383838",x"383838",x"383838",x"707070",x"b4b4b4",x"8c8c8c",x"7c7c7c",x"646464",x"646464",x"7c7c7c",x"9c9c00",x"383838",x"545454",x"545454",x"646464",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",
x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"545454",x"8c8c8c",x"dcdcdc",x"d0d0d0",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"9c9c00",x"707070",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"7c7c7c",x"8c8c8c",x"9c9c00",x"8c8c8c",x"545454",x"383838",x"202020",x"383838",x"484848",x"707070",x"a8a8a8",x"fcf420",x"fcf420",x"dcdcdc",x"dcdcdc",x"dcdcdc",x"d0d0d0",x"d0d0d0",x"dcdcdc",x"ccc400",x"706c00",x"383838",x"383838",x"545454",x"8c8c8c",x"707070",x"646464",x"646464",x"545454",x"484848",x"585400",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",
x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"545454",x"707070",x"a8a8a8",x"d0d0d0",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"989898",x"8c8c8c",x"646464",x"646464",x"545454",x"383838",x"202020",x"2c2c2c",x"383838",x"a8a8a8",x"fcf420",x"ccc400",x"9c9c00",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"9c9c00",x"707070",x"585400",x"202020",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",
x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"545454",x"484848",x"8c8c8c",x"d0d0d0",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"989898",x"707070",x"989898",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"848400",x"545454",x"545454",x"383838",x"202020",x"2c2c2c",x"484848",x"a8a8a8",x"ccc400",x"848400",x"7c7c7c",x"a8a8a8",x"8c8c8c",x"e4d800",x"e4d800",x"8c8c8c",x"9c9c00",x"545454",x"706c00",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",
x"545454",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"545454",x"484848",x"707070",x"c0c0c0",x"8c8c8c",x"a8a8a8",x"989898",x"ccc400",x"9c9c00",x"707070",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"706c00",x"545454",x"707070",x"484848",x"202020",x"2c2c2c",x"484848",x"a8a8a8",x"e4d800",x"848400",x"7c7c7c",x"8c8c8c",x"ccc400",x"e4d800",x"7c7c7c",x"8c8c8c",x"848400",x"545454",x"585400",x"383838",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",x"202020",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",
x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"2c2c2c",x"202020",x"545454",x"484848",x"c0c0c0",x"c0c0c0",x"848400",x"8c8c8c",x"9c9c00",x"848400",x"a8a8a8",x"707070",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"707070",x"646464",x"545454",x"545454",x"202020",x"202020",x"484848",x"e4d800",x"e4d800",x"7c7c7c",x"7c7c7c",x"a8a8a8",x"e4d800",x"e4d800",x"707070",x"8c8c8c",x"706c00",x"545454",x"383838",x"383838",x"484848",x"e4d800",x"b4ac00",x"b4ac00",x"646464",x"545454",x"484848",x"545454",x"7c7c7c",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",x"989898",
x"d0d0d0",x"ccc400",x"b4ac00",x"dcdcdc",x"dcdcdc",x"ccc400",x"9c9c00",x"707070",x"707070",x"383838",x"202020",x"545454",x"484848",x"8c8c8c",x"c0c0c0",x"706c00",x"646464",x"989898",x"646464",x"8c8c8c",x"707070",x"707070",x"a8a8a8",x"8c8c8c",x"707070",x"8c8c8c",x"707070",x"484848",x"202020",x"202020",x"484848",x"e4d800",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"9c9c00",x"706c00",x"646464",x"a8a8a8",x"8c8c8c",x"545454",x"383838",x"383838",x"383838",x"b4ac00",x"b4ac00",x"848400",x"646464",x"2c2c2c",x"484848",x"7c7c7c",x"c0c0c0",x"ccc400",x"ccc400",x"ccc400",x"dcdcdc",x"b4ac00",x"a8a8a8",x"a8a8a8",x"ccc400",x"ccc400",x"ccc400",x"dcdcdc",
x"ccc400",x"b4ac00",x"848400",x"b4ac00",x"b4ac00",x"9c9c00",x"706c00",x"545454",x"707070",x"383838",x"202020",x"545454",x"484848",x"707070",x"989898",x"646464",x"646464",x"8c8c8c",x"8c8c8c",x"707070",x"8c8c8c",x"545454",x"8c8c8c",x"707070",x"545454",x"707070",x"545454",x"484848",x"202020",x"202020",x"484848",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"e4d800",x"646464",x"646464",x"646464",x"545454",x"545454",x"545454",x"383838",x"202020",x"383838",x"9c9c00",x"848400",x"545454",x"646464",x"202020",x"484848",x"989898",x"ccc400",x"ccc400",x"ccc400",x"7c7c7c",x"e4d800",x"9c9c00",x"7c7c7c",x"a8a8a8",x"ccc400",x"9c9c00",x"848400",x"707070",
x"b4ac00",x"848400",x"a8a8a8",x"b4ac00",x"9c9c00",x"848400",x"706c00",x"545454",x"707070",x"383838",x"202020",x"484848",x"545454",x"484848",x"989898",x"989898",x"707070",x"8c8c8c",x"646464",x"707070",x"707070",x"707070",x"707070",x"545454",x"707070",x"545454",x"484848",x"2c2c2c",x"202020",x"202020",x"2c2c2c",x"a8a8a8",x"8c8c8c",x"707070",x"8c8c8c",x"707070",x"545454",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"202020",x"646464",x"9c9c00",x"848400",x"707070",x"545454",x"202020",x"484848",x"989898",x"ccc400",x"ccc400",x"7c7c7c",x"989898",x"9c9c00",x"9c9c00",x"7c7c7c",x"989898",x"ccc400",x"9c9c00",x"848400",x"707070",
x"848400",x"a8a8a8",x"8c8c8c",x"b4ac00",x"9c9c00",x"706c00",x"706c00",x"545454",x"545454",x"383838",x"202020",x"484848",x"545454",x"484848",x"646464",x"545454",x"545454",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"8c8c8c",x"707070",x"383838",x"383838",x"383838",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"646464",x"8c8c8c",x"848400",x"8c8c8c",x"545454",x"202020",x"484848",x"989898",x"a8a8a8",x"7c7c7c",x"8c8c8c",x"989898",x"9c9c00",x"7c7c7c",x"7c7c7c",x"a8a8a8",x"ccc400",x"9c9c00",x"848400",x"989898",
x"a8a8a8",x"8c8c8c",x"a8a8a8",x"b4ac00",x"706c00",x"545454",x"545454",x"8c8c8c",x"545454",x"383838",x"202020",x"484848",x"545454",x"484848",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"383838",x"545454",x"383838",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"545454",x"202020",x"484848",x"8c8c8c",x"a8a8a8",x"989898",x"a8a8a8",x"989898",x"a8a8a8",x"7c7c7c",x"a8a8a8",x"7c7c7c",x"a8a8a8",x"9c9c00",x"706c00",x"707070",
x"8c8c8c",x"a8a8a8",x"7c7c7c",x"7c7c7c",x"545454",x"707070",x"8c8c8c",x"707070",x"545454",x"383838",x"202020",x"383838",x"545454",x"545454",x"484848",x"383838",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"8c8c8c",x"8c8c8c",x"989898",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"7c7c7c",x"545454",x"2c2c2c",x"383838",x"646464",x"c0c0c0",x"dcdcdc",x"a8a8a8",x"c0c0c0",x"646464",x"202020",x"484848",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"e4d800",x"989898",x"8c8c8c",x"a8a8a8",x"989898",x"a8a8a8",x"a8a8a8",x"7c7c7c",x"7c7c7c",x"989898",
x"8c8c8c",x"ccc400",x"9c9c00",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"646464",x"484848",x"383838",x"202020",x"383838",x"8c8c8c",x"ccc400",x"ccc400",x"b4ac00",x"9c9c00",x"8c8c8c",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"383838",x"484848",x"646464",x"9c9c00",x"ccc400",x"ccc400",x"ccc400",x"b4ac00",x"d0d0d0",x"ececec",x"ececec",x"ececec",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"b4ac00",x"9c9c00",x"848400",x"202020",x"383838",x"7c7c7c",x"dcdcdc",x"c0c0c0",x"dcdcdc",x"a8a8a8",x"707070",x"202020",x"484848",x"7c7c7c",x"989898",x"a8a8a8",x"989898",x"8c8c8c",x"a8a8a8",x"989898",x"e4d800",x"989898",x"7c7c7c",x"a8a8a8",x"989898",x"a8a8a8",
x"8c8c8c",x"9c9c00",x"848400",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"646464",x"484848",x"383838",x"202020",x"383838",x"ccc400",x"b4ac00",x"b4ac00",x"9c9c00",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"383838",x"545454",x"484848",x"9c9c00",x"ccc400",x"b4ac00",x"707070",x"989898",x"a8a8a8",x"a8a8a8",x"989898",x"a8a8a8",x"989898",x"9c9c00",x"7c7c7c",x"9c9c00",x"848400",x"9c9c00",x"848400",x"706c00",x"202020",x"383838",x"8c8c8c",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"c0c0c0",x"e4d800",x"202020",x"484848",x"e4d800",x"a8a8a8",x"989898",x"a8a8a8",x"989898",x"e4d800",x"e4d800",x"7c7c7c",x"a8a8a8",x"989898",x"989898",x"a8a8a8",x"989898",
x"989898",x"848400",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"707070",x"545454",x"383838",x"383838",x"202020",x"383838",x"b4ac00",x"9c9c00",x"848400",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"202020",x"545454",x"484848",x"989898",x"ececec",x"989898",x"989898",x"9c9c00",x"989898",x"ccc400",x"a8a8a8",x"989898",x"989898",x"7c7c7c",x"a8a8a8",x"848400",x"7c7c7c",x"9c9c00",x"706c00",x"585400",x"202020",x"383838",x"8c8c8c",x"e4d800",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"9c9c00",x"202020",x"484848",x"9c9c00",x"585400",x"707070",x"646464",x"e4d800",x"b4ac00",x"848400",x"706c00",x"585400",x"707070",x"707070",x"545454",x"707070",
x"646464",x"646464",x"646464",x"646464",x"646464",x"545454",x"484848",x"383838",x"383838",x"383838",x"202020",x"383838",x"b4ac00",x"848400",x"646464",x"646464",x"989898",x"848400",x"9c9c00",x"706c00",x"646464",x"202020",x"484848",x"484848",x"989898",x"ececec",x"e4d800",x"a8a8a8",x"989898",x"ccc400",x"848400",x"989898",x"ccc400",x"ccc400",x"a8a8a8",x"989898",x"848400",x"a8a8a8",x"848400",x"646464",x"585400",x"202020",x"383838",x"8c8c8c",x"b4ac00",x"707070",x"8c8c8c",x"a8a8a8",x"706c00",x"202020",x"484848",x"585400",x"383838",x"383838",x"484848",x"585400",x"585400",x"585400",x"585400",x"484848",x"484848",x"545454",x"545454",x"545454",
x"545454",x"484848",x"484848",x"383838",x"383838",x"383838",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"383838",x"b4ac00",x"848400",x"646464",x"989898",x"989898",x"7c7c7c",x"848400",x"706c00",x"646464",x"202020",x"484848",x"484848",x"989898",x"ececec",x"ccc400",x"a8a8a8",x"ccc400",x"9c9c00",x"7c7c7c",x"989898",x"ccc400",x"848400",x"989898",x"a8a8a8",x"989898",x"989898",x"7c7c7c",x"646464",x"404000",x"202020",x"383838",x"8c8c8c",x"707070",x"8c8c8c",x"a8a8a8",x"dcdcdc",x"585400",x"202020",x"484848",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"383838",x"383838",x"484848",
x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"484848",x"484848",x"484848",x"ececec",x"646464",x"989898",x"a8a8a8",x"848400",x"8c8c8c",x"848400",x"706c00",x"646464",x"202020",x"383838",x"484848",x"989898",x"ececec",x"b4ac00",x"989898",x"ccc400",x"706c00",x"7c7c7c",x"a8a8a8",x"989898",x"a8a8a8",x"989898",x"7c7c7c",x"b4ac00",x"848400",x"7c7c7c",x"646464",x"404000",x"202020",x"383838",x"e4d800",x"ececec",x"a8a8a8",x"dcdcdc",x"a8a8a8",x"545454",x"202020",x"484848",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",
x"484848",x"646464",x"646464",x"707070",x"8c8c8c",x"989898",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"484848",x"202020",x"ececec",x"989898",x"989898",x"a8a8a8",x"848400",x"8c8c8c",x"646464",x"7c7c7c",x"646464",x"404000",x"202020",x"484848",x"989898",x"ececec",x"b4ac00",x"a8a8a8",x"9c9c00",x"706c00",x"7c7c7c",x"989898",x"7c7c7c",x"989898",x"a8a8a8",x"989898",x"b4ac00",x"848400",x"7c7c7c",x"545454",x"404000",x"202020",x"383838",x"b4ac00",x"ececec",x"c0c0c0",x"c0c0c0",x"a8a8a8",x"545454",x"202020",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",
x"646464",x"8c8c8c",x"b4b4b4",x"b4ac00",x"b4ac00",x"8c8c8c",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"646464",x"202020",x"ececec",x"a8a8a8",x"d0d0d0",x"8c8c8c",x"706c00",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"646464",x"404000",x"202020",x"484848",x"989898",x"ececec",x"a8a8a8",x"ccc400",x"9c9c00",x"706c00",x"7c7c7c",x"989898",x"a8a8a8",x"a8a8a8",x"989898",x"a8a8a8",x"b4ac00",x"848400",x"8c8c8c",x"545454",x"404000",x"202020",x"706c00",x"9c9c00",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"b4ac00",x"545454",x"202020",x"484848",x"706c00",x"9c9c00",x"9c9c00",x"9c9c00",x"b4ac00",x"b4ac00",x"848400",x"848400",x"484848",x"484848",x"484848",x"484848",x"545454",
x"646464",x"b4b4b4",x"b4ac00",x"b4ac00",x"848400",x"646464",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"484848",x"202020",x"ececec",x"a8a8a8",x"989898",x"a8a8a8",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"8c8c8c",x"646464",x"404000",x"202020",x"484848",x"7c7c7c",x"989898",x"ccc400",x"9c9c00",x"706c00",x"707070",x"7c7c7c",x"a8a8a8",x"989898",x"989898",x"7c7c7c",x"989898",x"b4ac00",x"848400",x"646464",x"545454",x"404000",x"202020",x"383838",x"9c9c00",x"dcdcdc",x"dcdcdc",x"b4ac00",x"9c9c00",x"545454",x"202020",x"484848",x"707070",x"9c9c00",x"706c00",x"9c9c00",x"9c9c00",x"9c9c00",x"b4ac00",x"b4ac00",x"b4ac00",x"848400",x"989898",x"383838",x"545454",
x"646464",x"b4ac00",x"9c9c00",x"848400",x"646464",x"8c8c8c",x"a8a8a8",x"b4ac00",x"b4ac00",x"707070",x"646464",x"202020",x"ececec",x"d0d0d0",x"a8a8a8",x"989898",x"a8a8a8",x"848400",x"8c8c8c",x"a8a8a8",x"646464",x"404000",x"202020",x"383838",x"545454",x"989898",x"9c9c00",x"706c00",x"7c7c7c",x"7c7c7c",x"8c8c8c",x"989898",x"a8a8a8",x"7c7c7c",x"989898",x"7c7c7c",x"b4ac00",x"848400",x"707070",x"484848",x"383838",x"202020",x"383838",x"9c9c00",x"dcdcdc",x"a8a8a8",x"b4ac00",x"706c00",x"545454",x"202020",x"484848",x"989898",x"707070",x"707070",x"9c9c00",x"9c9c00",x"848400",x"848400",x"706c00",x"706c00",x"706c00",x"7c7c7c",x"383838",x"545454",
x"646464",x"b4ac00",x"9c9c00",x"707070",x"707070",x"a8a8a8",x"707070",x"b4ac00",x"848400",x"707070",x"646464",x"202020",x"ececec",x"989898",x"8c8c8c",x"989898",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"646464",x"404000",x"202020",x"2c2c2c",x"545454",x"a8a8a8",x"ececec",x"a8a8a8",x"ccc400",x"ccc400",x"9c9c00",x"8c8c8c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"b4ac00",x"848400",x"646464",x"484848",x"2c2c2c",x"202020",x"706c00",x"8c8c8c",x"d0d0d0",x"c0c0c0",x"b4ac00",x"585400",x"545454",x"202020",x"484848",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"9c9c00",x"706c00",x"707070",x"707070",x"585400",x"646464",x"707070",x"646464",x"383838",x"484848",
x"646464",x"707070",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"707070",x"8c8c8c",x"b4ac00",x"706c00",x"707070",x"545454",x"202020",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"989898",x"a8a8a8",x"a8a8a8",x"7c7c7c",x"646464",x"404000",x"202020",x"2c2c2c",x"545454",x"8c8c8c",x"ececec",x"c0c0c0",x"ccc400",x"848400",x"706c00",x"7c7c7c",x"989898",x"989898",x"8c8c8c",x"a8a8a8",x"9c9c00",x"848400",x"646464",x"484848",x"202020",x"202020",x"9c9c00",x"8c8c8c",x"d0d0d0",x"a8a8a8",x"848400",x"706c00",x"404000",x"202020",x"484848",x"d0d0d0",x"a8a8a8",x"8c8c8c",x"9c9c00",x"706c00",x"8c8c8c",x"7c7c7c",x"989898",x"646464",x"989898",x"646464",x"383838",x"484848",
x"646464",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"a8a8a8",x"b4ac00",x"9c9c00",x"706c00",x"707070",x"545454",x"202020",x"dcdcdc",x"c0c0c0",x"7c7c7c",x"989898",x"ccc400",x"b4ac00",x"7c7c7c",x"8c8c8c",x"646464",x"404000",x"202020",x"202020",x"484848",x"707070",x"d0d0d0",x"c0c0c0",x"848400",x"706c00",x"646464",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"989898",x"b4ac00",x"9c9c00",x"646464",x"646464",x"383838",x"202020",x"202020",x"484848",x"8c8c8c",x"d0d0d0",x"8c8c8c",x"706c00",x"585400",x"404000",x"202020",x"484848",x"c0c0c0",x"a8a8a8",x"a8a8a8",x"9c9c00",x"706c00",x"7c7c7c",x"8c8c8c",x"989898",x"989898",x"a8a8a8",x"545454",x"383838",x"484848",
x"646464",x"dcdcdc",x"989898",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"848400",x"706c00",x"706c00",x"707070",x"545454",x"202020",x"c0c0c0",x"dcdcdc",x"8c8c8c",x"989898",x"b4ac00",x"848400",x"8c8c8c",x"a8a8a8",x"646464",x"404000",x"404000",x"202020",x"484848",x"545454",x"b4b4b4",x"dcdcdc",x"706c00",x"646464",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"848400",x"646464",x"646464",x"646464",x"707070",x"383838",x"202020",x"383838",x"484848",x"7c7c7c",x"a8a8a8",x"7c7c7c",x"706c00",x"404000",x"585400",x"383838",x"484848",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"9c9c00",x"848400",x"707070",x"989898",x"7c7c7c",x"707070",x"989898",x"545454",x"383838",x"383838",
x"646464",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"989898",x"706c00",x"706c00",x"707070",x"707070",x"545454",x"202020",x"b4b4b4",x"dcdcdc",x"7c7c7c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"646464",x"404000",x"404000",x"202020",x"383838",x"545454",x"8c8c8c",x"c0c0c0",x"989898",x"7c7c7c",x"7c7c7c",x"707070",x"707070",x"707070",x"646464",x"646464",x"707070",x"707070",x"545454",x"383838",x"202020",x"383838",x"484848",x"545454",x"383838",x"383838",x"585400",x"585400",x"383838",x"383838",x"484848",x"707070",x"545454",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"383838",x"383838",
x"646464",x"dcdcdc",x"b4b4b4",x"8c8c8c",x"b4ac00",x"848400",x"8c8c8c",x"707070",x"8c8c8c",x"989898",x"545454",x"202020",x"989898",x"dcdcdc",x"a8a8a8",x"7c7c7c",x"a8a8a8",x"a8a8a8",x"7c7c7c",x"8c8c8c",x"646464",x"545454",x"404000",x"202020",x"383838",x"545454",x"484848",x"8c8c8c",x"8c8c8c",x"707070",x"707070",x"545454",x"545454",x"484848",x"202020",x"404000",x"484848",x"545454",x"484848",x"202020",x"202020",x"383838",x"484848",x"545454",x"484848",x"484848",x"383838",x"383838",x"383838",x"484848",x"484848",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"383838",
x"646464",x"dcdcdc",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"989898",x"8c8c8c",x"b4ac00",x"9c9c00",x"707070",x"545454",x"202020",x"7c7c7c",x"dcdcdc",x"989898",x"989898",x"a8a8a8",x"8c8c8c",x"646464",x"8c8c8c",x"7c7c7c",x"545454",x"404000",x"202020",x"2c2c2c",x"484848",x"484848",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",
x"646464",x"dcdcdc",x"b4ac00",x"b4ac00",x"989898",x"8c8c8c",x"b4ac00",x"9c9c00",x"848400",x"707070",x"545454",x"202020",x"545454",x"ececec",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"7c7c7c",x"545454",x"585400",x"202020",x"2c2c2c",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"484848",x"484848",x"545454",x"545454",x"646464",x"646464",x"646464",x"707070",x"707070",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"848400",x"848400",x"848400",x"848400",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"383838",x"545454",
x"646464",x"b4ac00",x"b4ac00",x"848400",x"a8a8a8",x"989898",x"9c9c00",x"706c00",x"706c00",x"646464",x"545454",x"202020",x"484848",x"ececec",x"989898",x"8c8c8c",x"9c9c00",x"7c7c7c",x"8c8c8c",x"7c7c7c",x"7c7c7c",x"545454",x"585400",x"202020",x"2c2c2c",x"383838",x"646464",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"848400",x"7c7c7c",x"7c7c7c",x"8c8c8c",x"989898",x"989898",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"b4b4b4",x"b4b4b4",x"ccc400",x"ccc400",x"ccc400",x"b4ac00",x"848400",x"c0c0c0",x"c0c0c0",x"e4d800",x"b4ac00",x"c0c0c0",x"ccc400",x"b4ac00",x"848400",x"c0c0c0",x"7c7c7c",x"383838",x"545454",
x"646464",x"b4ac00",x"848400",x"7c7c7c",x"989898",x"989898",x"8c8c8c",x"706c00",x"706c00",x"646464",x"202020",x"2c2c2c",x"484848",x"ececec",x"a8a8a8",x"8c8c8c",x"848400",x"646464",x"a8a8a8",x"8c8c8c",x"646464",x"545454",x"585400",x"202020",x"202020",x"383838",x"706c00",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"9c9c00",x"a8a8a8",x"c0c0c0",x"a8a8a8",x"c0c0c0",x"989898",x"c0c0c0",x"a8a8a8",x"c0c0c0",x"c0c0c0",x"c0c0c0",x"ccc400",x"b4ac00",x"848400",x"848400",x"848400",x"b4b4b4",x"b4b4b4",x"e4d800",x"b4ac00",x"c0c0c0",x"c0c0c0",x"b4ac00",x"b4ac00",x"b4ac00",x"848400",x"646464",x"2c2c2c",x"484848",
x"646464",x"b4ac00",x"848400",x"7c7c7c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"545454",x"202020",x"2c2c2c",x"484848",x"ececec",x"8c8c8c",x"a8a8a8",x"646464",x"646464",x"8c8c8c",x"8c8c8c",x"646464",x"545454",x"585400",x"202020",x"202020",x"383838",x"706c00",x"ccc400",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"848400",x"a8a8a8",x"c0c0c0",x"a8a8a8",x"a8a8a8",x"c0c0c0",x"ccc400",x"9c9c00",x"989898",x"a8a8a8",x"989898",x"b4ac00",x"848400",x"a8a8a8",x"989898",x"ccc400",x"ccc400",x"b4ac00",x"7c7c7c",x"8c8c8c",x"c0c0c0",x"b4ac00",x"9c9c00",x"b4ac00",x"848400",x"7c7c7c",x"545454",x"2c2c2c",x"484848",
x"646464",x"b4ac00",x"848400",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"545454",x"202020",x"383838",x"484848",x"dcdcdc",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"646464",x"545454",x"404000",x"202020",x"202020",x"383838",x"2c2c2c",x"b4ac00",x"b4ac00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"848400",x"706c00",x"8c8c8c",x"c0c0c0",x"a8a8a8",x"a8a8a8",x"9c9c00",x"9c9c00",x"a8a8a8",x"a8a8a8",x"989898",x"c0c0c0",x"989898",x"a8a8a8",x"ccc400",x"b4ac00",x"b4ac00",x"7c7c7c",x"8c8c8c",x"989898",x"a8a8a8",x"707070",x"707070",x"b4ac00",x"707070",x"707070",x"545454",x"2c2c2c",x"383838",
x"484848",x"848400",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"646464",x"545454",x"202020",x"383838",x"484848",x"d0d0d0",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"646464",x"545454",x"383838",x"202020",x"202020",x"383838",x"2c2c2c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"9c9c00",x"848400",x"9c9c00",x"848400",x"848400",x"706c00",x"706c00",x"707070",x"a8a8a8",x"c0c0c0",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"989898",x"c0c0c0",x"989898",x"989898",x"a8a8a8",x"ccc400",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"989898",x"a8a8a8",x"a8a8a8",x"989898",x"8c8c8c",x"8c8c8c",x"b4ac00",x"707070",x"707070",x"545454",x"2c2c2c",x"383838",
x"484848",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"646464",x"545454",x"545454",x"202020",x"2c2c2c",x"383838",x"484848",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"646464",x"545454",x"383838",x"202020",x"202020",x"383838",x"2c2c2c",x"c0c0c0",x"dcdcdc",x"c0c0c0",x"9c9c00",x"706c00",x"706c00",x"706c00",x"706c00",x"707070",x"707070",x"8c8c8c",x"a8a8a8",x"c0c0c0",x"8c8c8c",x"b4b4b4",x"8c8c8c",x"989898",x"989898",x"ccc400",x"ccc400",x"989898",x"8c8c8c",x"7c7c7c",x"707070",x"8c8c8c",x"8c8c8c",x"e4d800",x"b4ac00",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"b4ac00",x"707070",x"707070",x"545454",x"2c2c2c",x"383838",
x"484848",x"7c7c7c",x"7c7c7c",x"707070",x"646464",x"545454",x"545454",x"545454",x"545454",x"202020",x"2c2c2c",x"383838",x"484848",x"989898",x"989898",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"707070",x"646464",x"545454",x"383838",x"202020",x"202020",x"383838",x"2c2c2c",x"b4b4b4",x"dcdcdc",x"d0d0d0",x"848400",x"707070",x"707070",x"707070",x"707070",x"7c7c7c",x"989898",x"8c8c8c",x"9c9c00",x"a8a8a8",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"b4b4b4",x"ccc400",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"989898",x"b4b4b4",x"b4ac00",x"848400",x"a8a8a8",x"989898",x"989898",x"707070",x"707070",x"707070",x"545454",x"202020",x"383838",
x"484848",x"383838",x"202020",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"202020",x"383838",x"484848",x"484848",x"7c7c7c",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"545454",x"545454",x"383838",x"202020",x"202020",x"383838",x"2c2c2c",x"a8a8a8",x"dcdcdc",x"d0d0d0",x"707070",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"b4ac00",x"b4ac00",x"848400",x"b4b4b4",x"8c8c8c",x"8c8c8c",x"b4b4b4",x"989898",x"a8a8a8",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"b4ac00",x"a8a8a8",x"b4ac00",x"a8a8a8",x"989898",x"b4b4b4",x"b4ac00",x"848400",x"989898",x"a8a8a8",x"a8a8a8",x"989898",x"b4ac00",x"b4ac00",x"707070",x"545454",x"202020",x"383838",
x"545454",x"545454",x"545454",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"2c2c2c",x"202020",x"2c2c2c",x"383838",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"8c8c8c",x"d0d0d0",x"b4b4b4",x"8c8c8c",x"b4b4b4",x"989898",x"b4b4b4",x"b4ac00",x"b4ac00",x"706c00",x"8c8c8c",x"b4b4b4",x"8c8c8c",x"b4b4b4",x"989898",x"8c8c8c",x"8c8c8c",x"e4d800",x"b4ac00",x"706c00",x"989898",x"a8a8a8",x"c0c0c0",x"989898",x"a8a8a8",x"989898",x"989898",x"a8a8a8",x"989898",x"8c8c8c",x"8c8c8c",x"b4b4b4",x"7c7c7c",x"707070",x"545454",x"202020",x"383838",
x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"484848",x"383838",x"383838",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"8c8c8c",x"989898",x"707070",x"707070",x"707070",x"707070",x"707070",x"848400",x"706c00",x"706c00",x"8c8c8c",x"a8a8a8",x"707070",x"7c7c7c",x"8c8c8c",x"b4b4b4",x"e4d800",x"b4ac00",x"706c00",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"989898",x"8c8c8c",x"8c8c8c",x"b4b4b4",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"ccc400",x"989898",x"8c8c8c",x"989898",x"707070",x"545454",x"202020",x"383838",
x"484848",x"7c7c7c",x"a8a8a8",x"ccc400",x"ccc400",x"ccc400",x"9c9c00",x"8c8c8c",x"646464",x"484848",x"484848",x"545454",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"545454",x"484848",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"545454",x"707070",x"707070",x"7c7c7c",x"8c8c8c",x"b4ac00",x"b4b4b4",x"706c00",x"706c00",x"7c7c7c",x"7c7c7c",x"707070",x"646464",x"7c7c7c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"7c7c7c",x"7c7c7c",x"b4b4b4",x"7c7c7c",x"646464",x"7c7c7c",x"7c7c7c",x"646464",x"545454",x"202020",x"383838",
x"484848",x"a8a8a8",x"ccc400",x"e4d800",x"ccc400",x"ccc400",x"ccc400",x"ccc400",x"b4ac00",x"9c9c00",x"a8a8a8",x"8c8c8c",x"707070",x"646464",x"545454",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"545454",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"484848",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"545454",x"202020",x"2c2c2c",x"383838",
x"484848",x"a8a8a8",x"ccc400",x"e4d800",x"b4ac00",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"989898",x"a8a8a8",x"c0c0c0",x"b4ac00",x"e4d800",x"e4d800",x"ccc400",x"ccc400",x"ccc400",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"b4ac00",x"848400",x"707070",x"7c7c7c",x"707070",x"646464",x"646464",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"383838",x"484848",
x"484848",x"a8a8a8",x"c0c0c0",x"989898",x"b4ac00",x"989898",x"c0c0c0",x"c0c0c0",x"b4b4b4",x"c0c0c0",x"b4b4b4",x"c0c0c0",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"9c9c00",x"848400",x"8c8c8c",x"8c8c8c",x"c0c0c0",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"484848",x"545454",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"383838",x"484848",x"484848",
x"484848",x"a8a8a8",x"c0c0c0",x"c0c0c0",x"989898",x"c0c0c0",x"b4b4b4",x"a8a8a8",x"a8a8a8",x"989898",x"c0c0c0",x"a8a8a8",x"b4b4b4",x"c0c0c0",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"848400",x"848400",x"848400",x"8c8c8c",x"989898",x"c0c0c0",x"dcdcdc",x"e4d800",x"e4d800",x"8c8c8c",x"c0c0c0",x"7c7c7c",x"383838",x"484848",x"545454",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"484848",x"484848",x"545454",
x"484848",x"a8a8a8",x"b4b4b4",x"d0d0d0",x"c0c0c0",x"b4b4b4",x"c0c0c0",x"e4d800",x"b4ac00",x"848400",x"b4b4b4",x"b4b4b4",x"d0d0d0",x"a8a8a8",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"ccc400",x"9c9c00",x"989898",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"8c8c8c",x"b4b4b4",x"a8a8a8",x"8c8c8c",x"e4d800",x"848400",x"8c8c8c",x"7c7c7c",x"646464",x"202020",x"383838",x"545454",x"484848",x"848400",x"b4ac00",x"b4ac00",x"b4ac00",x"646464",x"484848",x"484848",x"484848",x"545454",x"545454",x"545454",x"706c00",x"b4ac00",x"9c9c00",x"848400",x"706c00",x"706c00",x"585400",x"484848",x"484848",x"484848",x"484848",x"484848",x"545454",x"545454",x"545454",x"545454",
x"484848",x"a8a8a8",x"c0c0c0",x"c0c0c0",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"b4ac00",x"848400",x"585400",x"c0c0c0",x"a8a8a8",x"c0c0c0",x"d0d0d0",x"a8a8a8",x"a8a8a8",x"a8a8a8",x"d0d0d0",x"c0c0c0",x"c0c0c0",x"a8a8a8",x"c0c0c0",x"a8a8a8",x"d0d0d0",x"a8a8a8",x"7c7c7c",x"a8a8a8",x"d0d0d0",x"a8a8a8",x"8c8c8c",x"8c8c8c",x"646464",x"545454",x"202020",x"383838",x"484848",x"484848",x"b4ac00",x"848400",x"848400",x"848400",x"646464",x"dcdcdc",x"dcdcdc",x"b4b4b4",x"545454",x"545454",x"9c9c00",x"ccc400",x"ccc400",x"ccc400",x"9c9c00",x"7c7c7c",x"ccc400",x"a8a8a8",x"a8a8a8",x"d0d0d0",x"ccc400",x"b4b4b4",x"989898",x"7c7c7c",x"484848",x"484848",x"545454",
x"484848",x"a8a8a8",x"8c8c8c",x"707070",x"646464",x"646464",x"646464",x"848400",x"585400",x"707070",x"7c7c7c",x"707070",x"646464",x"707070",x"7c7c7c",x"707070",x"646464",x"646464",x"646464",x"707070",x"7c7c7c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"7c7c7c",x"646464",x"646464",x"646464",x"646464",x"646464",x"646464",x"545454",x"545454",x"383838",x"202020",x"383838",x"484848",x"646464",x"848400",x"848400",x"706c00",x"646464",x"b4b4b4",x"b4b4b4",x"b4b4b4",x"646464",x"545454",x"8c8c8c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"7c7c7c",x"a8a8a8",x"a8a8a8",x"8c8c8c",x"ccc400",x"9c9c00",x"707070",x"a8a8a8",x"dcdcdc",x"989898",x"202020",x"545454",
x"484848",x"8c8c8c",x"646464",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"202020",x"2c2c2c",x"484848",x"b4b4b4",x"848400",x"706c00",x"646464",x"989898",x"646464",x"989898",x"8c8c8c",x"646464",x"484848",x"8c8c8c",x"8c8c8c",x"a8a8a8",x"8c8c8c",x"a8a8a8",x"ccc400",x"ccc400",x"a8a8a8",x"a8a8a8",x"9c9c00",x"848400",x"707070",x"8c8c8c",x"a8a8a8",x"545454",x"202020",x"545454",
x"484848",x"383838",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"2c2c2c",x"484848",x"383838",x"404000",x"585400",x"545454",x"646464",x"646464",x"646464",x"646464",x"646464",x"484848",x"646464",x"646464",x"989898",x"a8a8a8",x"ccc400",x"ccc400",x"9c9c00",x"7c7c7c",x"a8a8a8",x"848400",x"707070",x"707070",x"8c8c8c",x"8c8c8c",x"545454",x"202020",x"545454",
x"545454",x"484848",x"383838",x"383838",x"383838",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"2c2c2c",x"383838",x"484848",x"404000",x"404000",x"383838",x"202020",x"202020",x"202020",x"202020",x"202020",x"383838",x"484848",x"545454",x"545454",x"706c00",x"585400",x"545454",x"545454",x"545454",x"706c00",x"585400",x"545454",x"545454",x"545454",x"545454",x"545454",x"202020",x"545454",
x"545454",x"545454",x"545454",x"545454",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"484848",x"484848",x"484848",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"484848",x"484848",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"202020",x"545454",
x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838",x"383838"



);

signal tex_data_sig : unsigned (7 downto 0) ;

begin 

--process (clk)
--
--begin
--
--if (rising_edge(clk)) then
--	side_out <= side_in;
--	bool_out <= bool_in;
--	texNum_out <= texNum_in;
--	texNum2_out <= texNum2_in;
--	
--end if;


--end process; 

process(tex_addr)
begin
	
	tex_data <=ROM(to_integer(tex_addr));
	
end process;

end rtl;