// nios_interface_0.v

// Generated using ACDS version 12.1 177 at 2013.04.28.00:50:59

`timescale 1 ps / 1 ps
module nios_interface_0 (
		input  wire         clk,           //          clock.clk
		input  wire         reset_n,       //               .reset_n
		input  wire         read,          // avalon_slave_0.read
		input  wire         write,         //               .write
		input  wire         chipselect,    //               .chipselect
		input  wire [4:0]   address,       //               .address
		input  wire [31:0]  writedata,     //               .writedata
		output wire [31:0]  readdata,      //               .readdata
		input  wire [31:0]  hardware_data, //    conduit_end.export
		output wire         ctrl,          //               .export
		output wire [255:0] nios_data      //               .export
	);

	niosInterface nios_interface_0_inst (
		.clk           (clk),           //          clock.clk
		.reset_n       (reset_n),       //               .reset_n
		.read          (read),          // avalon_slave_0.read
		.write         (write),         //               .write
		.chipselect    (chipselect),    //               .chipselect
		.address       (address),       //               .address
		.writedata     (writedata),     //               .writedata
		.readdata      (readdata),      //               .readdata
		.hardware_data (hardware_data), //    conduit_end.export
		.ctrl          (ctrl),          //               .export
		.nios_data     (nios_data)      //               .export
	);

endmodule
