��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ��>�(Ŗ�XV���=�<4����>c���t����֪� ��?��A������.�.��G� ��{~�޻9zZ��/a���<A�Q%�W��F�8�"�uRȸX*�V@��L���uZ�5t.yѤ���lN�t(�����.�}��
�9r��w�R��}����\qDu��d?e��r��y�ޣ�y�$�5Kȕ�7O�Q�g�������R�ɧو*B���UR<��5;_n���ݵ9,�!��*�w����#��t�0ߠDS���g�.Q#�S���b#it�`B{3�����)o��Ǉ>��~���ƉK�D�%	�30�1	@Y��G|@��ņ(��W;J���.�v�+&@�f�{�=�R��S�	e\-%�>*1~�C��1�E�yRN���QNN����"=�j
] �H��-Rh-��� �M-x����jSa�xKU�k`�.b�j����:��}H��Ѯ�#����uR�G�}�
��se)jڣȪx��:��Bi�B.Ě,��x9��@U��~�����Nl���;m��H��˓8���M��&,"�z*���$�4(L>}�5�~y�*�
,,��g��J��N��=VR�f�٪���ǔx�MĒ#��Դ� ��m_�Ef���:t� ?sؐ#�̲�]�RY�,�Xw���B0+�-$�=H�I���桶6'
q/�z�����+�P�����/��U�Jb�v؃o��m�}>%3�PCU�=�}O�z0�C�^��K��!�^��p�(��5�%r1~B�5C����z������.���m�TDM�"�XK�zz'-��|���%o�rͰ���2�ս�ּ[4�Q���kUj0S*��-��Em��M��&��"�:�8�����v�K�wc���e���9 �*��\	2#U)R�t���v@�k��,I�,F�uU|�V_��j�1����̛��%�p��s���<: A�t�$���zv�X���Z�`�Ki�/�%;��� L���2�.���Z�� �w�r��Y�)�[��~7�0|�6�3�y#ȵ��@	�pj���Ʒn��G��?�Q�F�yEԀ��"W�n����?j�v�#���hd�ʻ���l��Н�OFHZz��<�V�:$Xt;@���x>4`�ƐB�r�l��q���T���]������N4=i9p��$�B�#����-o���+�V������+��5Xxt�J43�κ�裂d'U�f��T���D�ֿ���S�ũ��Z?�k�taz�M�-�vQr�?�/���'���)��p���a��?��~S������U:�s��mJ��7��1l8?%�&T����������vDZ �4�=��bE,�gd;�b܂x(�9���'���s�x���gj�6�⽶]!���u<����)�)��(�ˀ��3�s[�|1y"%���V%�7�f�D��jB��TQ?��_�f�lA�[m����WW7uq���T�xg�wi���H~�UWu��P[�d��4ꙣ`��[�Ԇ���:��Q�$�b<ŝ���3t���c�y������X6�yx�N2~����H�UQ�L�OǶ�������)H������/�vޙU�	Zr�G@�Th�>����@�1�w2�c�����	�ť��w�{���ŗ��Ҳ�bL�Yl~x�-���(�@+յ���	^�늍���j_����diΡ����? -H�������?b3)ڻ�<�hJ�_G��?�����f �g�%Z���������:�i�nG��`�Ry������:;!�<������m�Ä)u�2��y�2�}���*-{j�*�R����39m�ۜo�:�1������y�@/��g#� ��o�cN��p�(J`��}n"z�S�G�k[�O�����B�
�l�6�� �c0�����C)`S�GUԞ��)�y���M�2��{���A)�[���Kf[3�R ��yƆ`�SYM%�8:'���4ܓ�G�0���HY��c��&I��W�_�bԋx��"�I�j>��]�j����m_��y=1�u7�=�	<��5�}�Ĩ�o�D��U�~��fD;�TP3��P��B��d�/q#HB5��d���r{'Kj5N����f!ж�+�5_k{��ظ�мA X�l���]p$ҽ�J!�Z���v#�YAM���c�O�!U�Vt�+���:�S$7,��ziq&��7��C&�m߈X\ߎ������֩D�����0�?_@ �Gl�Z�	uDe(��*�1[�B�� �>Z���6�=��6��J�J+������-���b{�O$-�������竎�mqYk�5T���Ə>�Z��#��� 1ҏ�3[��+���c�Y9$u�ڪ2�±���H�+��!|����7D%k�o���!&\��ԉ�/�{Go�m���9*u+U���G�o�؛������a�`ֶn+El����`0L���SX�5�2�&<"��Zvץ'(u*ib1 �LC�~����?j���"'<�����Y�}H܆�`���h��f/����^(��*�����A���H���Ί����	=8_���//�@�p�_�H�s>?���lHj·{]�P�Í��ok	�&��p�a��� �^�?5��EE1aXA_�8p/��㖑_��N��!1��b=X0�z��P�}���ϋ�y�"G-%l�ξ��^���7�{��`��@5=�r���"�WC%�V�N��).��$T!<�q?E�f���9��������k��=�F���r�g��~���;�8�k퇣��>�"͎2D�YO_�I*�w�V^f	Y�o���s���QSϳ�;��.q)604`�s<r�6voh&����QO�^�qxL�����u��n}��% ��-p�����	QJ<R�(���������]!��fT�T��7�ь�ň�^�%<�lS�m�#-Y����0q�]�.ŷn�����@��叉~6'���N��["ݯ�SՑ�ޚS4��| �yFJȴ��D��Y�dR�*�H� R^]���4�x��BP��2`4^�9\N�At�3�=7���ғ��x���g�t��P��:�Sb~�.A"�1X����� C�ߧY�Q��ߣ���%�d���� g�e���n�� %���� V���K:�d�0�%� CJ��~&:��q�c(4
�@M� �6�� T�X�����,3=�뎞�)`�5�
K��?�,uX8=�AW�W��`S�
E�y�-4;j<	��s��k�����6@��1�°_�>�^�Ǥ,yg�
���fͯc�ys�|K)�b��믍���@lgP�I�)',H�;��*NYu�.%��:5`��i@~5���S��˥&`e@M�����?7�N�e��2�p�q���tHrf��#@�4N���#6�_p�,��V��M�{�c�		���+Qc;,eY6I=i�Y�'pa҉��1�6CEQ����_��ht��f�8�����_/�H��gU��icp͌�(
ҏ�hрd�^LKg���)��C�;�{��y��b8��00���KK�*([�g�,�]��T�U�:`M�p"�g��}H���:���ġ�g<L��=9q�����L�|��x/�K�p�>fUP��� ��8�U��q�_���LB���z#����S�u-~ū�fd4	�%J�T�ɖ5^b��V���G:�8�`��N���[��z(�3�q��>2�E�I� Hjjs}�U���Z5T%́�jpҮ� [,��r nR$`R�Y#QB��E;?�G������\��W���\�����!TFk�(8� T򻓯p�pn��
)���0WJ�c�Z �٢�.��iP�/�:���	��gl�!�BoƤNd/m[�u�/K�.���eƷ���~Ta	;*�@ER֧�*o:���ŮDX7wZT�w��l�{��G������3,Hwө�.� I�p�^]����
[�5�)�K-.LG2ץ���?�bl���U�oub���69�������D�;��e��UZ��K�&�F�!f�u�T�E�Lm����SGp	��~���͘޲u��ī��F�����x�8P'��R�OR	�
�;�7eP*+D���'��ɤ��D��k����ۣΘ��@�m����(sd7P��7X&v4<_x��jJ\.� ��ό�0�Tr>4�;�����mm���A�V�#h[�%7�����ӰR�`�����A����Q�1@�"T�~m��(�=�u�y�w����@�#!C�w'��Tc��Y?����fڌ8�Je ��\�=�h�*@$r�Vfq� �*i���Z�d�٭�����JpKe�D$��b�<���Wz����K��OF��t�Z�I��Ơ~�֫@`To[Vc+=5�n�ݨ��5��*��(lԢ&�<��q�������� Z�K�7��gr#[���}2��1�뱮��#�,�dS�n����A�^GR%e'u2R%�ik?|�x\���O%�~�	���5'A=�c��n��Q�w-�>��<�͚U�.l]C�H�TZ%��	������k38��jVe�ɴ�����nH���y��+H�Yo�U�s�V�/ڂ�	����'Z���C�>K�@.�GK�t�j�u�$B����E�"��n���X+�.��]2���I;��?���q���D�8�+��\��#Y`?����V65�k[���SQ�mE�$��t i˟�M�Wiy�w�P> �4{� �Rc����6A/Á .3,�~�]!���'a�T��ݖ����m�:j�r�_���f�7�̱����D��-n�g��b9,r�P����!�.k���ݙ��/�W7�?;���^��v8>T Q�N_A��}�γ��1{p}��||�-~;2nYk��a�C��x*�5h��҂q5V��wU��*2_�Y��%0���?o�Hz�B㢺C�EÈ(k%Q�P��{	`�M�&�1"���x=�V�qɖ��l�Bs5��k[ꂾA��H�)��O��=D����C�����DI���f��ۜf�A.��3(�b (-��mYh)�B.h�2
�5�u� �M�ޡ��|H�S�BW�4!�V�H�����!� 4�u�k���wY.o
�+���yy/���1k��³C��d$qf%�D �w������4���˂�V�"���Ȃ�&"$�ia���k�.%�ٲ^b;��SxW�5���J�h\z[D�@W��j��_��.^��|�ڊTؔ��1�1��)sF{��� �"����,H��|�aJ�,[�㑯�R$��f����2<�@k���9�$�ϥ�݋99�0���g��,ap8h/x�]��k��iZ���쒩��<2��	���� ���'2x��Ż�D!]����@���+Oq�g T_Ɓw�uKX�En���^Ci�$[\L�e��I��ń�t�({�Y�ko�0<"i.f#�A��9��d�Me�H����2���@�eş�-�4�h�d�"�:�j����������e�����s
n����ey�Q`�m: ��_/	�]�>#@��'I�tOLr�W+��\�0���\ ��W&���&�p�Ci�,b��u�{�|̬�l��&'WC���ˠOe�鶀����T�Wڢ�̦�2J`R_M[Je$6��}����If�HD�;&�q��4�?�����o��8Z�����X]�Kj�nϗi�V�BM�C�����������k�2�i���X�C���H�B��4bK��u���W��ώ��^��~��p����gr_��;�F7_��M�\
�i�B�ȵb_�%l�/g�#�)�jj=w��XK�
�H��Da?1]��'����x�Fê�m�Б6X��d-�`(�rF.��-�Xϙ�Mܫ�j��"ko�����4�������c��6H������Z���8�bL���Cl�Y{
���~�3?_�Ё,8�H��jp��6��P\���wFv@N�`!���!�3�Yy�G��#�9k�;p�Ts����� $�	�jYΝ��Rp׈gR���
���`�jU���c���c��xN�#]�<�2�%^=hP���{K�[غ�$�y*
L B���s�`�$�'�_�����8ɾǶ^KY$	N�B���Eb������@J��}v�UD1Lb6j��p�,,�.{�m+)R��.�sf�V�`�`N=��f�<d���bh�I� U�0'�������#*(�ܣE��%Bn�`t*B���OȌ�z$�}߉չ���sim �P����D~�m���vgѤ���	Jj�_��R	�w�d��=�[3����� R�n������h�\T�Xx���5�%�it_��;�+���zσ����hTѰ-����﯂i�60$}��W��`%^�t}��6ƿ�[���$�0f��iETn�N�b�^n�MarY&��M�[�@�KD\���_��(�������d��(HŎ��!r�u�����ϩ�wD�j�S:�����^�Q��O:�Ë]�bt|��@Yn�}Ѭ��y*�iiR�qn�n��~A[��\MrT�+�}�:୆_�B��
/l:��#�u�����j0��@��c�F%bT�Q04�Y�":�Q�"��x[uٸ�W���Č������UO7���7�L���8Ѡ��$������&2Rpd��=�s"��K��ӷjAe�&z��\4��`�ҥԍ��*�6�I`ʋ��rꈒ���jy�d�6!����`��b�˺����4-�)�2e���EG'P�c��W��̡��L;�,���`S���q���{�!����=Q�"ں�����c�t�f%A�q�c^+��tԴ�����{�#P���7d���ԛ��bp�x�f@ևP��/;�o�ȵ�Gy��V���qsWF�����_�1k�'�b]�x�6)fp:M���R��j,9P!��P��OcA��ż'���'Sмc����uA�r��R��O`���	,i�N�N�n+0�m�gKOCc	^��D���uc-��j��d��|�/����+f^g_�v���$w�ie������u7 �r=Y+^#q�f �1�E�]� ��,A$�׻����Mm�LJ���j�Wr$,۾�Z�͢T�k�zY�h��-�P�
��vъ��`�v1����Uv+�4�h�x�1$���|WZu���m䳜E%H2§6[T<+��'�4�{�ꟽ�c"�v%�<�N6���h@�r��N�Ҝs�Wڷ|���m~0����RwO��p��ؐ�$C� #X�����P�H���#z7翛TB�@�h�m*����˫w�?��i7���{j�+9۷�՛֌R��a��t����/-P��歑��:�<^sp]���+BT#L��G�o�j��f7|���ߜ5�Č�
�.qh0>�QҊ�6��8ގ��ek�d]�nO��v7���*���}���s6UnumA��V9･[���wR������e�z�FD Z�6��sL�@Ȼ���+H3������^�3�h�[C����ߕ�@���y��y@���)O@=ƭ-���FE����i&Ao1���)��μ �/XjxpY��V�p�ʲ�Ң�y�H=�Y,	I���%GeT����g dh	��T�3�5[1��h���z<����~&}�>x��S��\hr1���5��X��]�)M{��d�d��R\����S.!N.u�K��Ƭ|o1�*@��D���s4t��]8]��Ȩa���1��w�9Imzo�wg@���w�:�G���H��څ�6b�	���������X��
���q�����Kݦ:(1�Ș�K�IJ�h�9E�e�F�8
�Y�BV�D 7�P2Op��P@w%a�bhL�*���P�-��D�����|3h\9N��R��C�~@���>��>'�J�f�h����6M	�ǐ_!�~?A�D�5�̸Ϧ2����[D����}7�IPW�茫�/�k%oS�����`b��}�!�zẅ=N��%��c���UyO�)I��@%_׆^*��b�]��wnrN�'��qD�p��7X�e�5��n�cǯ�o��%�pU�}��:�J(�͘K4��W¦,`������9r�.��p�/5���UP��O�6˃�����&�ƥ�Ǡ֬����&�A�_�x��R� � kot��@�M�|����3�O�SP�~���Jw�.E� w���t%%��u��:��{�a�⊟�����t�ܐ'��.Wc0I5�C�av��0����g;�ć���Q���W\vJ� s�&zj�E
]������΋����R���h�������q�N*+�7��1����(�s���$�ZŅ�X���(�g�Z���pF�]iWS���r�-�K.(Ch���yحUU�f�R�,QLsg@���J�raN��R>Y7b]f�|�����چ�+,�.AmR1���S���������JB��b-Uۆ>���ݒaz��+�����43!����S��+���|x����� V�v�2Ȳ���!��;�ZL���b3\�[ њq�o١�a~���?�ֻ�Gd��:Y�"�� 1,(�|0�Vo��ZBH��;UCY  �x�314�{`�ML)��{2�"���r޼�M=����R$�YC
����\saztW��H��%Wj�i�Ouw`'U��;L�x������a%������#�1�%�ϲ`�*�e/k���Ɓh��� K-[��,dA2��n��)�Kʄ�x�k��q*�����盽^C"��KA�c���^9�ѳ�����R3��t��k�ȚA'dY�%��OS��Y�,���G���RT J��Vb��{L2�zC�1�v���֜�"�7�6رj���b�sh,��_3r��������b(Rhų���8P�ϝ��HH��:�OZـ��N�d��:�bOq�0��=��됎>T�iR`_z��c���D>d�5%�V���-�����U2�Z��֪��&@���<&,h��$f�Q������?,P��o�k/�Ap9kF	7l�̔o�{.��%%�P�Ɔ����{�y�{����zm�_�V"Y�T�M��7��,q��X*�F�Y|��B� �h����cV���ܳ�i���3SI�fVw>��69c���P�I3ۍx_Q�:"݂NUZ��}�k��bY�I�n��p�u���b���}�4�,�gM��o�('���b|���7�T���<\Z����V�o�����ʏ��D�nt�ц����/��
z�8_��&��%"�L`�RX�jv���.�댯�!�*��"�Rq��r�vy� ;�"��ɽ���ޮ�s#�kCv�����o_�D�B/]��;\&�S����n�ѣ[�|o�&p��L�Q�'y�2�骪e(@25%�
D�8p�ޞV>�/no��&��᩟���}I����dɽ�ױul��)�p���*�������pf��n1��V�^f�6���ke��Tv��qi��TQI�BO���݊�4�d�2�h�$F���4o�;�n�"q�isz̪B�h� �)W��Mx���&o���B����l���7��j�I >4�Z�w��h�t�'�Yx�#�p��Wܱ|g�6�E����D��=�x�-���a�)�r.Q��#���#ژ6�@Sd�:�B�+f=�M�܇U�t�m;��\�,1��6�̬���J��Ʌ�*5:���R�Fzt	y�n�L"*�u[���񱿦��Rշ$��?)��5A�`z����ؠ��0MVG���:��m �K������f�b]�pH�5'�N���K{<�| �;9@�͡��U��`��\n�
Mj=񤷪f�j�F�w6ڤ��8�,��s�}k �Ð��9=�n�P���^��սmg_�I��]F��	@��X%���<'���M���,xoK�Up y̙�3֎��1��=m�s��*�?�ֽI���!�:p�7��NI�X�b]?�П��G�TsO��g��� 7'�/�b��®e���7�E*�V�B��O�)*��
�,��kjғ��K��Dӻ�\����>�B�Qc��k��Uw_�pBҽ\��@/t�ޖ��K}ԭ<d1���jqDZ�U,ى�u�Y��n(��:�6b�Bl�7�r�SL@��9�-���	X��z�9%�z����AN���0��4�r��U�����ݭ����qA��;Gtς {#q'N=z�\��ڢ<�'���"M�������L�1��0��v@Hē3��Os������|���4����-��ڋ��FϚ�;���.N�B�w���Em#�_Q���i��(S����ә|=�Ƽ��F#Uj�+���u���قY���m¥���_N�#���p���gkr�qS��l"�`���z�����y��u^k�Q_��	��0 �,���m�t�]I5����s���X�IidfO,�o�Z3�����9���]��b���s4�o�@s{���}�;�.�1%��WVC�A�9վ��K�}���%�����(��)�!Ey�� �-����"r����x�n�8�<IT,��.(���t�	�CO�yʟ×�`v�+� ��5����JA���G���Q�Rf�K�N��Rɺ�Y�~#bɹ�&ɻ���Kz_�����yt�2�q��?�$ ?�����2���v����a9�XL�T-�4sQ`����x+�B����Nl#�����(c�*��
���*`z:D�*�锶	�18���n��5�oT��6�����G�����?�K�\�27F�p�����ԧ����"���U`%�$��m���C'�m��'��dܩ\ީ g�#F���1_���	I_�8T�`�����u��ЅбW#���+e����҆���%CK�izq����]����lحJx$o�psp
��+����, [p�itEs�J>X$�ɸ������>��?�o����i�3���ä�%�,�}�#��=�=?�N)��0�,1~�}�#�YNi#X"R#��������"�Y�z& �Wf� 7���۫d'-)q�QZ܆r�1��؁�'����.�͋�Hn�x��<�Ը����aMh�1�a)#ut)�����I�>!�����Ȫ�E�Hg��~�
��/��^yv�uk�Y�	z9��$}'w��uc�se�!��b�VA� �U�ܦ��),3k�i>����8Y�6G����9��c�Lf��t��3�tY��8����l3������Y���췜�f'4S�g�[AȌ�n�o�\��˿k�	. 2�_��1)fS��0���j�r��7�i�v_���@��j�0S%��)���ī9Fi���KYC�S
Cp�VK�3�͋jn��g����)U�D@������2u	��ͧ6܀/֐�{MCՍ�r\տd/[iM�0y4���0U����B�����֔�ɖG���aU�m�ZCP\�:�$<�mS�)?a�H�;10I��$x���Bg�sX���&���J5�S1RU�sY#?_*�XY>Z���`�T����F�İ��r�w9ρWm�3�t%ߋf�9op��Ԝ�Ƀ+8�����������.5 ?hf)� ���U��..�w�r�m0MlN0�cɃ�8��YD1�(ɗns?	z�ݮ8������E�U���tA痲���!Cu�?�@g��	hg&�]4_MT�Bx��	�%J_��xO|5J\�^�r�'L��K{��`&�޻=��Y� ���ܺ���n��,� �uN%3S���t��"D�f}�5觳~)67T�Za���Uc�o�'#ЅzO�^E�uW���F�o��s���}}��ac��Q�D�r��O�_�5�<H�>srcăW�G�0¹����|U�C����Jx���9O/��MtޣZ>E��֟�\
>B0-�]�a8q	2�@�G��V����m���4���3
��$o����V���*��C�{�9=П�A��ft\C�?�����7��_
��ǉ0�F�N�R*�Sic�KJԟ�P��������
N�(�]�����29�� m�=�:7��=��!���$��H���m�����-��	\6+*Vj#C����xa��,[�����܄crҒlPUEM���NQ�+HY�:���v҂S��+��ë[�	�{���R�`��7ݛqH
���U`
�i@a�z����
9`�1�Ǒm;��
@�,sB�lK��P4hLF�Jf�3�W�A��}5;G������\�����5��y��^�\����` ȸS����v���Mc]~o5;�Pж�����iQ��my@�$�-Dpp�����X@L��)&�p��J�#u�#^�/;�՞�/���iU��Q�D�e.i?��P�A����'sM|�u<�eY�	Z�֯iej�4�w���@s���_�~	�:ъ�o��*���Ԟ�4����a?�Cg)E4U���Y͑���]ޘ.�s�1B�qc-��
��Mr�54���È�LZ,�;q�/���V���P����@�J!�˦�~��~�$z���u�]'L-L�5�^�M��!�{�A��n	�*ǫ�g:O�*��g0#�<��-K�}������S�t���p�+"u����m����[~)�ۈ�Y!��nM*kZ-B��n�\p��]b�N@�����lܘ�o0��(Z�F���u�G���υ�pd��/OR�,;�<���*���7�|�9I`�Jq�=i(� ��/��<�����~	��q�hN4�*�j�-���ϝ<���!�� �T��@H� Ih�ZD���I��NH�b����4�m��#�b��#_��Ԟ����7���էȸv����M�Rg/C!5@�R�� ��@��z����iIfd2y����6\5?!7Z���>aiI�4�t�I%�3O��.ysK~}�P�E����|�A�nv{<z�x�΀O�%T��������L���nƆb�e�>9������X�������E%��-�F��x@����t3�Rb�U7V�ЏUE?,�д.�w,w��ܳ?#A>�w���ۯ_�Iu��e0�Q���+����&�'ʯ����(M2H����5��(v����<�`����BN�o���A�d����=M%m��kߤ��|��V%d�®�s~B�<V���t?�˼-��G�e�0y;�sL�7 _u10��d�~�n�E��C���pT����e��ֈR��^�� )��k���'e��@�↺��5j�K�o��G��ݟ���)(���<�/n���b���%�X0��h �t��l�����l���peH��E�^�r~p��d}J�ֲy��}	�C�s�vQ�t��R���goL����:�(�w�4 ʷ�(ʑ`�h?��܏�vP���'�NȽ����MB�L�����()��ʁ� RE!��lV05��>,!��"H�����~*�0�c�����@�����8���_q�~�ii��)�J������-�-i��� 
���2a,� ��}Nō�#�$-Y�9!M>0^[���$�.O�v�S��$���cB[>���4�����,�[xu�V'���q�Qq|V��Ӗ��l�f���h���eha�D۶ܛ#[�"QN��K��&t�m�-Ԓ̧B���9��%_O���f�RA�@f;�}���c,�+Qc #��p�A��o�kh�:���O�#v�E�b����C��`J�d��U�Z�����m��y7�����Jo��6���D�yF�����,�_[�s�U��N�~����]�J]��U�k=��=ܱH���%r�aP��<ۡڤ��&�a�[��?	���P�5�
e|�wn��(D^�i	�h�#��	�n��>������UOQ�w\x�R�a�Q@�2�&���vbS�>�P{Y�Wem����3b�9��=�w��K ��ͽO�� 5NQ��Ix@kk,��� nBcgV9��^�dq%qv�Vwm�� ���jct*�\����c��-��^_�]h���ƁS�>�Ҡ�@��~�.�ӌ�x-iȎ5���lb���ӵy�^�ǀ�-����M��J{����\!~"(�p��-�C�C����YO�i|���/$���_]��?(,�}���婫oC�#a/�M�K_ds�>X��b��x���V����A�鿍	9�#K{���4sb���6P�F)�83�����Q��_�ߌ�#�����:���.�b��M7%-%���t��˱�@D�+�Q:��s���?4�|��9�!E�jjp���%�U�WY�%��ߏ}�	�T��G��<s,YH���?�D*Bֆ��8�޹��4��wAS�CP-�:Ti�I ��H�F?�ڛ�3�`�d�Mp8�YK>����z�i�X����ZU�r�^���h�m�z��N@���@=Ֆ�bC]H�8%���� ��1�n4�������[�0�M����Ҽ��|}�e���k�3�<�?�Q�
��w�aL�^���}�[vȨ+S@�W/���lLA�%q�?�Rh�g뙯���כA�@��ޚj[�o~�5�Q�'ͤ��c���� y�ط��p��˧c�[�M"��L�p�Rj�\�����I��ȸ��A��iဟg��" �W{�
[o��b̑`�
:!b�uQ����Y���B����R�Y�f���s�A*"�+�G�b��֜�s�����}B�SAg������E<��i����+)�@�����JZc1i�F�
�v��� �IS�}�D
�2Nت9���$.��1�P������s<��p*�FI�����դ޹OT��T�UU���+=����UY����6��Ms�qB�e&��;�Fq��~��o�G�0����C+
�WW�س���+XĪZ��=~ox\$��m>�У���\v����z_$�mRg�n������>?d�g�C&��3[H��t,zά�䬹��Tq)�����~*GN�4>��J��.W>�� ��a�Vwt�X���d�|�&�/P�f�: ��~(�y���c0���U��pG��l���j�p�^���Qv�ǲ� V+W�5j�٭�"�X�g�����X�6���=BA
*a�Y�<i�ƶ�ѳ�-�`}��T
ih��Ѱ�<Y=.�+x�ԠA�S��'��=B!X"��Ic�2��Z���hT19�dM*=T����Y�_��
KcQ�J��YY
����״B�����k��h�N����*���xY��~Yr����^�ӉǼ�\�=g��M�v��5n�Ԥ�i~C*������V� �ZU8^wp�(���"��|��.CWM�f���� L��84;�P�$�/�i����wU�؂G��X<E�:6vH)Ъs�`N���{@]z�q:
t�D���ؖ�oH7�E ��m��K�kH �w4}��T_&��ȶ~J���Ά�m�S��`0�&�o�c��7�����{�}6�@����٥&U��dTGC#	���E�9�ی1��j���3�T�8��	��=���|��R%z�캋�533��g|r�6�:�JJ&�mh>a�
r:��V���9�gC�K����6T *�~թ�����Y7����%V��4h87*1v�U�Yߘ�o`g��X�x�L?n��4*��BN�y�|D�TAY0��<c\�-ʽҖ	�ho`R�,�V��]U@��^|M�����^��;ʖ|<��U�Z�]������ ѣ�c�*q/߶M���4k�z�h�H��$��0���6�0�5����,}���B!W�q����yF;�$y�̄3ec�d�zI����F��@8l��.g���n���VL(�����;��}������r�2:��`���ll�Tu2,dՖŦ�{UIZM�BW�}�G��U���}�'Α��o75�$d��k&�k��8o f�o�H�<3
W�]5�vgD�H�?~����2d����A3����>��n�Q_�A�Ð���ob���zO��3��A��S_�\���D�r{��ꅡ�s!�v�y�X:BLtF��S��&�B�ı�o�_."������B�6O�=�,eI��&��P��.�?t�y��+4��})��Ո�?��/!eKM�����������H���}��:b��yaB��������T\QS��>+�A��V���K��JxgIT+G�
�Tcg�"���-ՙ��̜mǪ��9V���sIRV/���bW��u+����V�@���E�K5Dь.r ��Wc�~�ʵm�@l�И�5����dc���j�����[�-�/�|ߴtj�qdO��B
��z�Yϻ,w������r>�v�v͈;%����S흵Wl������TT�ذ�p�ͨ:$���6ˢK��t�bL�FX�eTO�X�"_AsNn�(��N���&Dmg�V^c�o��s������|!anK�'4�7e�j;�zGM���YՁ2b�Ή���G�GϏJg�B=�
�_�w��b��LF뻗��/N�M�8V�CD��GR��%û��𒮲(��>�p̓Z��̃�
��}'e�3`����z
��u���gVz�Kţg�Ϝ�~��8�L���ۃ��[D��L��n���GΖr=���Kug�Dk��E��|�;@�hˤ7߭$�/�\g�'S�����g�*�h��C�	#"k�<m��2���|���.=E@8�J�T���N��6���@��ˊ�D�)O�G�B����e\���O�W~}�u�����@��]�>_J��n�D���T*MO��C��dI˂�����]n3�3�B�[��u5q�Л�.���#M��\J٪W0���(�2�o�}�1�KL���������#�k퍩����S�U������{�-�ğ8��d��z���� !m�D��O`{�6:�^� kEE�#��z|{�~��:?@����Q��h$v��UmOS�f���,�s��2��M(/�o���2��������󧂨���#<��V���1h�~��:�Vdu��@�;|ÑKч�����$xK�d�[wdE��Z@�������H�n^ڱ�@�߃~����"���R�Tf�j���;w ��@�Vrf9���a@D�q/C(��#i�՘���rI�*�����<;��� A�1�B86�$��l��d������:���	aӶ����Y�����QV�ޭeN����*Q ,�?��j���H�-p��nV�$�a���A������Q��(��`iE��C���z����j9�aS�-�N�Ȃ�8��
2k����Z���z��6��L{ۗz�xݗKU]@_���Z�M�P@��ߠ�L����F��i���c�M�
����k�GB�׮]&̓'͂uC�b��~vM�^�W�Dr��@Ty����� �)���n�Ϊؼ�.�H|E����C_�)(��֫��{sy":	>�K�3g���L p+54����J�!��mj+Z��$p0y#,��w4G4^~��Dpm�:Pzh3%9.�X@HKg�R�O���h�q����3�P��y�RŃ+ �roK��k�<�We���3�O�a�+��@\ީt B��a6�e\2���ˈ����܆�x�Ьj���]��;�_�]�{���89�N��2;EWt���Z�A��@�b���s~˲!'�]� ��j�8��W�ƈ	(W}�a�;LsW���<1% ��u�y)��q��Ц�=��4z�TgW�����p�>RƧP��%�u�����#���^�н#m-���`pk	|&�gVB�I�M)eP
��|�a��P�9��po�-1n���jW�{_��6�h̛w�K�U��*?z�N�w�F���΋~��%�m�h&e�����rӼ��*�P}�� -BN!i@#.���B�U�n��zn*�_t����=z��G�����X�u��h�li������+9Ѻ�z��4�����9�3���&��6��G�j�Ҏ��P˿-������A�}y��d)�F��D��4*���_O@v1/���	���>��)�ϥ�Pl�$a�;}ut�DQ��ܒ#��=��-)AϞ�,�7�sy���8�tJ$�7 �E��{!�ee�X��؎��NXT݉ ����'���`r�t��d>O�\A����
n�F���$��.���������-���Ib�ꬼ�jr�~əcW(�}uSu��l�`�W�J!��R�В1�*\�37��#Q����>x*	/��Z�7�)xdr�P�����ϫ����pz�������.@��s=%�ֹ=����N-�r��?Pq�M�(�0�R�`@\���w�:i��3[�h��J>-�Z��\�=���[�l�����/���ˣL����?�v>��M���Z�Ky�L��E@�H#��k�v�)0Sy�e�p5�p�q�t�JS
��T�&r@�H����F�����)�����V�]D��+(��'��e?�^0*6�YkP/(�ޞdp��untɉtZ������	��xǮ��|�6�|�W
31:9$R!�w�rG��m+��cu���VG��t`���G�wӿ�`U�x|B��[K
5��M�G	7���N 5K�0ֿ�0h*`	�k�H��.;a��"�5�Pc��1*5օn������%ڊ�kG�e��W���M���l�ۆl���3# p	2���m��~� ��2G�ܤ� �ѬI�n���΢��OL�F�
���4Q��8�x�Q,��>��[+Q���b��J�����{6��(��0�_�fB�%e6V�A^Z�
�w����5
���)|��h{3y��x��8�
ל�)�X؀��[��s��p=����OuU3�) B��=[)å��̘�|}p�v>/��W}YN��at]�<��i��y�E`y��$�	�' @�#-�8�=Ơ!7�Z��o�r�ƭ����֖]�`ˏ��[��=��x�C�EH�t��;�.C�AAٞ�!{�#N��.�ROӔ�2k��2���b���C�z9T����/�J�1L�+������m?v@��p����V������ko�(���������'Ȇ��B���1��u<�G�0���窜�Ic!F���ȬH�B�X_11�a}��]��gd��װ���L`�+�v�*���#3ݹ�%��������a�^QR���/iߗʏ��T��� ���@������^�� cÀ��-�7c����R^�܁��}&��4�]x^��O���wl��LDK�آ��9K�u�8)�a��3�C��%�ǜ[����g**mf�ϭ����%ԓ`��R(�E�����_���!R
���[oE�.�^�>H���P����sY	�>��K��F��:�z@�X9�(�?��iG��o��)�?f$��6ϣȂ#��*I}�c}��a��}���7��N��P���p�h�F��� @�W(6�4���]	�ɺ+x;"##���{�z|�q�ǂȆ��4:�b�N��_�#pg�U�]��4+'�Ufq� 叇����s�Ly�Dm\5d¡W�-6l� �(B��DbR�nnG��岒��n��2w��:aY�XiH,5���(I�m!�@��P��YC����M���^t�#6,+	��9T�%���S7���F�mJ�6Rf¤�7 B�����TN�ȶJex��{�H�g)NV�m{T�L��,"'L���}��$�����Q%ڌI�xut=���]�BWbP���9�,�*�����G�_dkvocՇ0Ǡ_�"�4�q,�݈��L���8��N��$%��6�d�ǧ�CzbO�͉��Y� �Z��!k}q�""�^���;c5�����aS�8F���g��`' ��T-B)9�5	��_�����~��h��RU���W������q�R��l���+eu���glN��]ų���;س��"��S�%c�;�
��?��Aw�Rv_��1}�Y�KT��q@���H�Z��Q� l]}�N��_�K!g��N����L��"��&�g� ��*�L#��y�K�m#��2�����m�<�h�B����Y~���p�W��&�M�D���j�1���i�z|xɼ�&���A,:K���,�O�/���{˿����](�깺�\̠�0
� �8�£������V��!�U��r"�Cշ�:�O�Ζ�R�ǂ %2��g[%K
񭗊�d���r��[�p�Ƴ�4SF��y��B�� ��2/�i�f�f���ϔa�h��ٺ�1�L��Z��ܼz�"������RU@��.��������_<]�n�Z�^�:;���XNFd�g?��t62<*�O ��j-tN:Jn���·BA��� <6�����h�&�`�/��n<VJ�֙�O�oK�X�t:@z�6��:�nd%]e>�f��� ��C�����Lu�����$��N-C��N��  �<0�&��0����{!�#:8C�[>�#C�3b^M�2W�WSQ� �J�q�LA͕���0��0ÿoO^�M(�LjLw�c��2�����	�o#9[1v�.���軶��
�X�Y�
������&�_O&���h��:�ޞ�j݄�=����cI���άd�T�����\��SP��cBc���*&�ށ�F�M�]�6�Ơ�7�x���_ʔA�⹝'ʓ��|X��e_SC���\=;_�-�^�T�b΅AS�����u�,�6�TC��
.��W�b���w�zB�����cgK|�_�s�� �D�e)���$�;��E��W��yLA��yf~s���9�X��U�4'>��/�]��w�^v�������a��J��V���"��<����E���Y��@���-��࠹�5���
��$��R��)����Y��c,�mV���`�m�	�<Uk������[�lRɥ�&%��.;+Ȧ$kl��?J{?/����W��g��Oj�S�Ro�z�mQ�7#�� �le���_�#��t��m��ZCp8é	q� {s݉�]Y=�fq?��/r�H��m���r=e*�&���q��#/�QG���W�I���� �.d��Z��x#��G%����c��ax��zAQ������L�d�BNb+�qutr�N��;Vɝ�j{�K���(/�أ���#���C��r���C~�%�����S�X=i�E��8��8�x�iwh!�1�1iƐeĤ���g��Kۻ��#ؾ}���SX�]5t�"���4��FD�$O������'gkC7���8x0l;E	&�4���k�z>�Z�_^�V&��(x�ha'ˊ��w/?�$
�����z� ^�Z�F�Ky�ࠦ?���zR�@�{`<�y_Ѽ�0��	��k9D�i�X��\���bg}gw�nQ?-)]�}h�D(�m�{�؀�A���~�w�(��ҏJp&���IX��O�E]t>���O�{�a�b�⤣��V�`�f���Y�	���Ì �*lql�yY��Ie_;c��$Ka*���:a\�j�e�L�q�e*�tq���:4�����m�bHoGL�R�J�J�ʒR\d31��+���g��lTfT���o�*�%�?�?@±�A3�V��1�`���֊�*B �I����X3����l��8��@-�5`����!�\�e�e���^��3O�e�ef�����bQ�V�x*tV%�z�*l��T��&�dB�}��Ox޳���l�紃�~��>V�c�,Z��CV�,[��2�˿��;ҥ5$C�..�4�e��y>�2Z�d_O�X	]�xX��vm6��8V]䳲 >,� ��C�t,
�갂v��^�&Ό�i-�u=��y�t���MHn�/�����9���ě���S�s�CWY�
0M�}�J�����&[����i��YE']�M����s�f�c��7Ǆ@���:��)�@ß���r���@٣kʽ���E��C�F���Ұ$b�`^3F̈p@Nk/\�T��� ��ǋmQM@9�ַ������Qqb��Ng��߬��}kmV@-h+����1����o��0��`�wT��+�bu�Q$ ֚�x��p�>b���M�y6 *�S�*�A�K#ӻE[|X���*�Fs���܄aU�9_��S'iE�5|��\���r��C�VYXB��)�Q�@4�t�Rb�@���*�2����:�UL-ci������3����M�z���N�~�|�9��h����*ڸ�����TH�Ǜ|��}ဨl��(/ƁX�ōk��D�"^�z�Pq>��J?b\���Y�o�O�x�"&��k�Yaܪ��[ȁ�VP�#$!	2d�/�8��JaQ$@�ҽ;y�d9d�<쯤B�l�g�����{a3݋������
��<��lgW�����6�؊��f�v����Kڑj��r�uȲ��R��Y��p�E]�������W�+��`�1�����ˑr�&��Xb�t�gc�/:�����.�,ʐ�rބ�p��B�mguY�ۦ[A��"6=�,�K�d�e��� t%H�������@����On�A��;�OJ���<�4��Y�b�Sf�N���jA� �� �G����e~ڨr�Y�.�Q`@�˭��A��Mgu�Sc\�w =�~	]����Y��x2�5�7��:���l}�0���2kĖz������=���;�]�̰�y�~�D����
��,M� :ۡ�z�)'�-�j�����\YlUo�����N9���8o���"LJ�H{/�V�� �Zs}�au�ˑX�i��[G���Ít�P�<<�OHT5�>�DNt�I�Ft�f��ғ������)�0%�j�>��98-�[�e�K��*}	n� ��K��ES�1�sz'�7Ǔ{���:�Df����p\���pGPX�n�</Lɝ_��o2z~����ڔ�����CI�[�i��õw�ڻ6j����p�C�?��oiF��6|:
�\�q�m��m�C�4Gk��Vܻ5��5�<Z~�c��K�Ss���J[rd����8�=|���TºRl_\��\^)�I\����"g���3�ixy��ٹ��V+JG�	!��Z�/ ��޸V��F��iƛJ�b���D/�K�H�y-��w!�%��փ��N$1F�;�f5�}�]`_�=��\� �t@���,��?��NzCF�XK����JN���/�q�T��S���pPs9��+���o��u��������v��P���@�&3����b���-�g=��F}s9�]ɭ�ƅ�Z�� 	���������b�޿��!�9�0J�P|���4=�^7��܋����1�����x��!Ğ��
�3U�q����Ohd !��S�5��z<k��Cp�ј����V"X0	�Vt�*��'�z�RY[.`M���H���<y	��*�,�%aȭ�@|�.�2%�����7��PN"y�BĆ���Z��RTO�Z�3��7E%,`�" ������T�ŘB*ѫT�6�K�g��6NW�W��c��ˆRꠌ��pٕt�G1S�i���x�Q�a���,�J���< �B��g���q�5'���:��c���x_�/�:K�h�-�@@�T*�}�����s{u�o ��E�
@ #d<a=�W��v����f�Y����!UH�Ԫ�c�,���xj��Ƹ��N�f]�����v�m�;���l��[oL�,�j���>Bp@����"	��V��~Q��ƃ�J��,eJw�z�2��L�{����gh(@��Z�sq+�S�Ӻ澠0�y��׷i\��/����[^�K��nr9oh��,>���%�!wn�.�J��i��\��{��}6oqϚ�bL�ڢFti� ����f�!%N��Yo�R�
�HX5���a!�Ѻ(��]���!׏��w�w�xY���@R��jŘx����t=�O�����I�F�����}��b�B�{�ť�W�Gq2��]����8	c�K��ҫ{D�Pʢ�w�w+�	Pӛ �&��FhI��{j4}5��� (�z
-ܘ&�efA� V�W��˳�'����-��܅���"���2%�5��D:z~1aSįX�����S`f�p��ߡ-��ԙ��Fd�Ё����-��҅�ۃ����\�ĥ���J� :[��︃�}j���C��7�º�5~�;V�u;��C���`/�P�d7'!Wi�����H����V���M7$�f��Xlx��5�H�W�qL���]����O���q�҉ �}$�����8�<��/U~N���5y��H�:_���I�����	����� �P�j^
��A�n<�=�	F?��<��5��:�=;\���J�o��.}���eFj�X/�DÖ�0bQ ������G�J�ѫ��_࿺���I:��Fm�W��ζ|z>��A���$�0��4[!�9s>���DQ���< �$m�hpR�E[����-��1M�d�lڶ��}�#w��L��D��rVL�)ٸ�e�lsZ�I�}�*b��G0+!�ϰfN� ,2뀫����Gc�9�ꭂK���X�8����D��������ڍ�7����/mq�	;�)X�0��<{26��f˽
�2�iN�$X�Z�˻��ԟ1MP�W��M�p�8|l�`]�(�������Is*_�ʛ%NO�`'�H�m ���i9����R*Y�Π
�=�rD,����w�!��&�15Wp4��e��O�NP@�>ƑQO$��؝K�b���Ց}^c�F�Bo����>"E�%�w��q�����QӔ����}�'�������eM@ȝ�;nF�	Vֶ��K� }��K��2�R���21e��M�0
��w,���RҘ>�!���
(L�7��be�6Θ,�!1�X�h�iK�U�����n�hJ7�e��u�uU�_�7	��b�J˲�L+�s~1
���b��ɸ��D�-Z?*+mn�GLJ�t^�4yZ奪�:���t�m�)35g�u0�ӄ�� �vEQw҉8!��$x�CZ���Dx�Y�E��|-W�t��%��:��r����>����ma���HKr�5	�T7����i^^1~4��[m�L��]���9W<��&�Ty�㻡��'HO�zT�5�Ur�r���>m�pN�Z�.��\�� ��\6��\h�o�x�ݱẾ��n��a��MHm�-��3�W�e�׋+%�����CQ:�e��~EF�4j�ӯ�̫�^�������M.�o���p���ܞ`>�+�l�亁'b�D��഻��?1�up���7$���`	ф�=
���ҞءQ˯�t|�B��G��� �$��W!�MX �4��^),���/ƞR�Е�8��qR�hNF��$��˼ ����A	Ū�ϟ8�b8?�{��I19cU���w�G�g��6<@w�f@�].@��{#\��\Њ��Y�����q���ߞ��BS�6��[�踊9����n%1"�-^AE����Wx+�,֚mC���4�'�$��Л��>�m�]m�o�� VN!Tz��d#��.�j_�&��4����_��Ll��u���N7*�}���E�����]<B�)�$'J\�8�'?#}Xĺz�^� 9�o)e�U���-1�@�� ��aYG��|s�i]������P/&B� VY�wd���ZCl�X+��b���=�"�'�L��/��k�W�q�(n��\hq�Q��px'=`=A��+:�"�+Ǭk�KtN�:�u9	�z�*��&���۾0�F��L���|�~b��"��(���>l��ا��̭jٮ��3�69��ٽG���&��N�4j}�#��p"���!q`OmK���=M�*��u4�������|+�R;v�1_E-@U�5�c�aof���o�&�3�4��cfd�h�O")��7ؤ����!+j�i'.�ǝ@�/���~�����t���q���!H~���u��j_��ʆZ�'[���{�}�'��v����$�L�u��
׹��h�t8 �;E��N���2��drG��iW��H���B�.�}3@'+���#�
-�cU�4ӿ�H�wp�-��pԫ�T��N�P_���w�$�W�c�#~'�Z��O��Kl$�ȏۻY�olsJ��/g"�h�����AG��18uY$#`IWF��`b_"�9�Ea�vx6l�(N�W�y�7��}��1�@9�Ќ8�n2��A��1q�M��z,�X z8[gn�<�*�D�0Y��
D@J�@���Nt�}�>B�>`� ��x��g�h���*�ua���o�?~0NyxԒ����)!��P��:���B�]�IM�����I`�=�EF��O�9���1q����h(w���o<�,�H ��Ɯ.%���;t����ێ�J2��j N�*�.Gr2��Ύ��:��u>��,�W�����������߁]��O�7�*���3���������N�"�pc6�����o��+H6�M��w�Ҵ[���TU�v;]6������ˣq��p�|v'��|f����bDDD�	���0�9�b����5Ŀ�P�n� L����n|�E��V�.0�Gp$��>|��kk�O�r����\/ov��Q��`����ym2�z/b�}fl�%��b�qs�����1���g��~6��r|P�v��N�~R�,]s���yQ��|_[����JO��dG�Ϳ��`���ˁ�E���Ls4S�;|�c�忧�v��NA.�;\%ueJ�v%�=H<&�\�D���a�>[��e��Il�Y�:�%i�n+��rT����e"Էp�"�8��%������S�����wM)����8�5�~��g�$Hɸ�SHMm��HÍL!���n�@�-�0��v�-�ba��Emĺج��`�re�_�ߟʅ݊|Of�2!O��ԫ�%�.v`٢�Ch����̍Y֘�vf�c:��4x�+��3�����/���>��� ����,�l���G�8p^{��$٨��s��:q���}R uٔ/��L����0

���?�|&_�ڼ��z�<�j�?Kj|�|��i �Je>�?�1���2�=��u�R�Ɖ,����#g_��������j;c�Iw���?{p��������T��U�aP�em��� q����aڿ�W�Opn'.����qptI�H+�9H:k�Z1<��
��lPȯ���L���q��;�A�_�?�/�񌯟��;4[MhH�8ظW����Ɣ�cY��	�l�G�9����$�V�wxɼ5���=�����L!;a����[��7�_���Kt��g�誎���5!E����U%�S'�� ]�����O���l}��#��Yo��l8��N�ry����q֗�V��ʩ7�~%�D�v;�,�f��AҒ���6�g�m[X��4�v�̫ת�]G���T�	ݼv�Y�'���U�Q���m�,���'��9��F_3Mߊ���41؜��0�횪=hr���q^$����n*'O+}��(��"׻L	f����^��5��"eq��V�.���u�X�F���7t�����h��]�s�#����jPW�@���,Mˡ�T�����M<�U�1����sC�ZB�Lͪ����v	�S�o"��Q!��z������n{�|�i#�
����V�տڔY����$�����r[ �������"D[�H[ ��/�h٫�{.[�48�	cM�G!_3�s��|�t������S�:N{F1\��_�m�e�}`,8~�w��>+�+Y-��G��	��pP
�S/p��61\�Y7��?� G�o�������F��n6��zE�ۼ�q�/j�;��T���Ke�o5�.Vgл���.��g�Y!D��F��w����N�1]C�IQ��0�=������)��뻗�n�>�* |zU�5��.7�<H��<W�}k�A�
�pj$��w�w��Sg'�.�'^~J�>&s�Me��a�VA����E��W�l/h_y�kT��Xk�7�]����ez�����N�#ti�ok�`1A�*�/�\\<���TTd~��yj̹��VB]_��Gf2���_�P��Yw�C>H�dC��k�q_�ݝ�CH��L\n�.(�b�r�hl0�$?l-T�	�b��]�I���E���׎�T���Ŷ�ě[&ܝb��6�8�O�f�J���P���0d�8����]��'�H��eHZ@g5ٳ��ڢ��_�;k��u�Tx��L���%�'š�����f����"�_�4�Oj�8�dB,m Ka�o7�	[�	x�_��7h
W[��R��'�xaﮆ��0��a$)�/����6����-N�j_�Z�aZ���� ��}��\���f��lp���>O`Q�4�q�c�K�����s��|���O8-N��O�c�����e<�HH_�7�=
dЙ��Oy�/܃��o�f��D�
�=M�y\�6�,����d��yG^����_eՕ[�̹�h���:�МR�5h��쮧 ��u�К;	�>Ɂ?��g_�tG�0���VjƬ�Y�νЮ�?����������	I�����|�X�cW���
��7���_�s�ހ�'_�Nb9�rbs�J\�}3��D�l��P�������{���Xy���`���Tv�a]� !N���VD�� ����Lx#�E�,��دq��0����?\K(����_�&��ר�<���?�u =DX'Jm~W��M��&'fR?,A��Y��d��v[q�U���C,��]�.�a����H�w�������
a��\wP�h{cs�Z;!D>B�p�aVG�k����Kr�դ�T��F;��
8����Ƽi� /Iy�(�gXQ 
��a*�`�Ȥ�����͒L�=�?�	;}A�A'C'yƻ�������C���xP��������Q�֞Mޯ��**j���65��o�<�L(j�,!C�"�D�{w�<�k�_u���, �
�T<|�/��h��ā$��X#�Sv-�|H�����ڽ���t
oh�
�*PT}��-�1R#em��-<A��Q��k>��F�B���w�)�@!`��:}`��ؠ5���(�x�DW���VEb*���=ڽ8���M���X2��O�yE�#��~ɟ�,S����c;�568	��-�
b�Ȁ�2aK�XJ-���ŤA~��x٫�W�+yT�W��u[���j{�=�%4�OǌP>�d4�̗����jU�pp9�X�p	U����A�e�CֿO�@a�`w��6��#�"�ۮ�V��&�s�E���[
�n�,G�g;���0��%�Iy!
n�(���h3}׵d�vn�d.���y��ʱ1�ch�Ed��5��������>ԙ�K�sx����:����_`g��y�ov���c"�i�&�f��!���"�����
��uF��S��v��%�dGCLS�:W��-`��f����,9��WSh��[L��_��+��&r�6���[��@��p=�RY��v��>�=�c�l�}N��@1ЀH��xN�ң-��<��
E���t|�Fʛ���&45�!O#���-��t>mvſ�RRR3�E�X��f#K��g\����A�	������BZ�(���۞���S��ډ�0B�鱥���QBtY�����'U���n�Z���ǚC��X�?�v.#b��Z;݁gs��`�1�nb��ͯ�X����o7O�Ӂ��~�#z�$�ϭ����8��_D�Q^����:޵�6��ZCOT1�03q�����Pɳ�s�f�3I�{	Vi����n{�@xя�j\��zfH]�h:� ����(L��p84���ͮ��4Z����N1�hB�h^�.z����mԝ#Inň��y�.�e�p��Չi�F��̵KZ)�:��4��Y��U�ur�@��9��:o����W��,Y�fI7Ĥ�?*�O/��ZwyT)K��Q�Q�<@1���p���m�=��dJŤ�sAD�*�<����"�~��q�����=	���d���n�)ԍ�����V>���o�
f�W󜃂~[N)�QF�_p�u�3�Z�k��=�b��A�F,Þ��R��[jt��U�g�7��K�7��⽄M�I�|Y\�dH����Q�}�c1i�@h�"ړ�n�X.�wX��z_��7DtV�s/�ݳI ?▥&��pYO-���A��D	&�h}�G�k`Czh2}��h,Q��/�ެ(9�@���1�Ť�'��{��c��'�z(�%è0>�'��՞-��h�vL�	�Z��5�&�7B�x�v}TU��0�5��/�͕$�����X���X�^��.ji7ǰ��5H�Г��}���4׌R����DI�ԕ�]���������ȧڮ�#Ca��xI�_����
�C�t�th�>�J��N�y�_����ߍԷb-vߍ.`�H�o���b�jGv�����}�Y����*��z�%F]�v@�q!�����C8�@פ�cn&PW��퐘r�^�Ӗ`�ju� o]-B���ܷE& +�e�tUq�Þ�c'
�&�	]S�iy��ɳ�Yr�]�ܤc�m�Ul�_C�� �=H����L��c3{��jƫ��KE�%�s��D\���g�n�u�n��6⁗�^|w[ұ�F�,@4�!2�)ZU�؈hyP+��?-�
I:��OY}V�>�Pm���
����uKb���*b�me$Lx�,,��Sq�1�zP���$�ٿ�?9.��Y�R[�c`׌2��j|�jff��MY?��{��l�_�,���[�^<=�������$�F�.w4������D�3a-�>4�����R�"��8-����n����p�H��M������-܎��4��KX�$__��L^�s��9�BKcIV��+%\N_�k>A9"�:绗z����[��8������b���ۙ;�S�"TP��P2X6sOA ��0��+8�P�O8}&�05u�:�� W�}>��-~A�z��j!���� �fl?�QU�
�M|.�ii9�_E4�?��C����{Ȋ$�*I��̳'��Y�x�`���563�y��R(o�}�b=$5��g�t�E�3�7ƞ�@�ƚ�ش-�y��� �.�>�_Bi��[�:�l�V�m���'-��ihd@��u���~چ���Z��i���y9ⵡ�ҥ}�.�Բ'��Pa\��H�vm\?��8���V�,�& 1�cI��IӒ�3n\�s"����4٫�]m��kÉ��:�w��������+S՜q�`��X�0|�-���"�<�ax���-��f������*Az2&x���p�#S��_è:M�(!2���Y�}?ML5���sŁeh-6��S�*4/�����'j#��\��uM�Y�0�����gP��[��pFX��Ä`bA�CZc^G���)AqK5sib�]s�l0�>��۸�(^p����}��f��ٰ����_K��j����bԙuw%���T�:�0(��۠5V\76�i�S�ى	��d�^P�_U��w�� fK:�:�xi���(mڑ��WۈKY��8��S��u,��չ�R�al�7�����%=`�]�p)u�s.c��ᙫ��D��L�'$Ӹv:�`�	�ԔV��@Ű���%֩^_kK��V-��q�PW۸�UC,H��+	@���	U��㶬��l.��Έq�͵��XmJ�d����� ^ς��~8�k�	!�O�҃-7��_Q�8�b���T*��(N����=�NAݴ�iN[��P?[�F����H6[�8z I+d�Ja�������w�A��|D6��P������ed���Y0��O��A#���>�p��Y�����a8UR��90�K���Q�4���&��ę�Վ�0�Yi��<��r����fb����0��=�q~��|�R`�3�G��
����[,�3.��4�A��AI8h��b�ß��}`��=^I#�v�Jہ �Q͇f�������~�X��ICN��L�u���ٟ��t�&����@��ӯ�%�z�]6�9I�5�s�z�$�m3)Knf�`K$�M[�0� ���k����
�}�,�sR(��@� �#��2�.,��}�#�~�������6dvC#f̵��'� ~��@B����-/�`�L��v���|V�D��g�;�,����s3qUq����ˣ*#����i�_i�2�����W�����k�Ľ�e1oo�� �]r�\�z�C��NO:��r��-`���D�d��D����h��)�չ�����s�����`��YZ�7y�M1$�m�m7yY�<���q�lw��h���qrʣ��=G�d����m�?���1 pw	�6�e��������~A���n����֛ީ��V�|���$D���Y�t4��
^J��+�5[@0�E�#�#e��5��+��u�P_�sX�L��.s��+rUlN[>��Iw�|=�{�����U"�+�����H��e��r�1"Ǎ�X�ȧ+�ԃz1�O�w����Z�h�4?49�>H��Jv�Z�v�¦�%�4��ˎ윷S,�(F9B#���.�3��Յ8G�ٔ�/w��첝���Gz�)�?k��fZ�q{��zW�^_~���H/�a;ű��5�-�BTl��Yt�1I{�M�(�".��Ҵ���F|����x�	tr���(�����>���/I�E��hd~NS�a�A�Z��oM_߃�e��g}�3�����&�
^P����5��d�t,%����Tr����63�ߒB_�O3>���1�ف��e4�QPy�s�ǳ!�8G=@u��أi�i�+�e3Q�8S3];�z��G`�>WǇ�V|�$�Y�/H���"B�i jXY*�^H�"gc�*��8�I:Q�ȏ��uc��V戆dX��BDR�M��@v��򩴫��7�_�lS?ĕ��z�H;}�x�q�]� �g< P�v�g���]$t�E.I�d�}.z�*�x8�����L������L؃�UP��n�F?$q�9K�N	�6�*g[���F�v~�-r2.R�Lkr�/i8���]E���6Z���&��]�Bh0�b(�^mԋ�*M9��+��3k��xP����H��r\Δ\��c�v��\����W��K@hz'�j��Ε�V� B��Ԅ���
��}�
~�+��7Нxz�3�>&�!L1�ް@�[:pga�i3�W�ջ��2Y�9Cf���n�æ����~V��a���7ƚ��UIL�+���9R>>�ˎ�œj#�k�T�@L<
����!��M9��H�T��(
�\��9�K�!P�6�Ƣ����jm�8�3�¶���f�HW�Ϛ���Ԕ;E&�ߋC�N��Y��w�2W�-~�7>�;o~=��C�̏�b�8��C��w s�*O?�����������1����M���&l�Z5��À�W��
5		[
'���0��]*$������)T�)�9��}�:�	�F&�9�`�.��6b�t^��y��.��Ә��*��<o�z֝���J/�c�"�{+�e/�(Ԓ�:��������G0>O��`��5��s"�J-��$C��*�E`��80�+�\8�g7��N#GK DpO����n_ 8]ꢚgyK�(@��ɻ�0��:�J�ab�V��F�V���������ͦq���	c�h������� i�yP���ä�dP=����̭�� ���;$��yV9��"�.R�|�1�ހ��n��2�8�����^mW�D��$��ckA��FG'�#vfb�)�Kf�2�8�,c���I�R���0b.3��%Ȋs��)��<S {(n�ۨIIhh�@I�ؔ�:���% �c�ѣl�p���~��΂�՛:��"�]���8��I�dF��Ek�8��iB %��s�mZ,3K3��Y��/��Bb\���,������(*�h�{�!?���b��tp{�c�<�0�Ax��C����ʁ�;�_,�f���U�����j����z!�Ԁ�9�U���20��#���$<��m�r�hrg���7��	�r�-��A�A�x�rv��v��K�`��::{w��<ß�`�g�'m�7lq�?%j�*�ݿ���S�+;�����V��ɭ����M�r�jlM���Y�uh�B��y�t������$O�i��+YS�+���@{޻��t
� �	��iU-��2�t�̷@��@���_�&�z^�y���=��Yϝ�s�/4|����m:+��Z�lh�]�_�����XU�)���!GC젰���+\��C&W�.�~������/�pO�唧����!�_�F�׿�*�CF���������As�_o��8��L^i[�p+ԀP^rOia��t���b)�� H�ۂ��~�	�v��k���ҝ�
68�xWN�9u:���jhh��Z�1� m����M-#�F	�5�,�.�L�XϯC�;.]w������>�L�=м��-���A�*�u��i��h�V��G�cfqjU�yu�}#��54��۲��sW<5M���z�0�<���*�扲�_��dg5����bAP���u+�e����:����_�zW3�$dV�ؑ�3�rt=�&��k�j�dqh��gOOBݙA�
��ߚ�)^�I�|&��Ԅ���o�v�>;�:r/�S0�S7��5<Y���Sĸ��I��9ݹk
'
����Hy�e~ z 1�s�G$�� �Æ�vtC���D��z����X$-E�g��;��u��o3�D����5�k�#->�'���G�,&�d��4`N��>�� �����G��E���*c� z��Q	���T��{�FsJW��H�=��Xr�kT��$4.����4��|P�Eݿ����̾zGVYQlb�J̻^��Y���}�Ou�#n͕�)�Ro)�9���E�[F�U��>J�[�՟�Ȭ�?# %0-:u�(<��5��.��u�����c/��
��4?-�\Y`��s��3\���*�yq���Vxߊv�m��gu��u����ϣ������ ���ץ4K�/�3]�H�� j[Έ�m�kᵏ,.�)�`��!�J>��&����vml�\��Êcu���K�,���N��K�ެ�_�ps�G��Oz���Vz\�3K��}=��c6���J��T�P�Ƀ��<�]&Ɖ�ĉ�M����W�	�QJ�|vl���̺P�#4C�`�^2� ����[� ����MO�V��l!~��dep�]-6��M+"mD�'�?���I�d����r�1��Ʉx�B½��Mj�H��nl &K�y���/�����t~��H[�����au�ŠM�.��<oS'�D۳�>���"���ќ�t��ur+	�$͡�c��.�	2�C٘��f�Ƒe��D�yA���(_�U�n
B���q)�X21�Ǘ<� y���c����2����#�g�R�a�CS��-�� r_� V
/��I���lOu�t�b�f#�0j��D���B�D��`/=����w���sײ�m���ϭ��󩁧�pT"H���	��1�����_�3�K�=��7Br��u�5��6��Y�u�p��D-5/g�tm��԰��f�� $���G6���4�G�^�5��[� �]-����*�xA�PS\w�o���r���f>1��لGPu�l�� �<������7��#�a�����N�y�P�Ě�1�w&e��܉���s��(;y�El67o�U'��4��pdr���>��_�*��^�H�U)��JI����+�p�]�%��[#p��_h%�	ӴG&�/)��F����p�\�V�;�U��x-ʉ�ʹ[�s~G͏^���L�� <6�$ޔ�w&l��L����W�`ඏ
6��ע�LyHD�ߛ���KM���
T�OB�(.���H�*nXG���{PN���Ě=�?^�,�H�h�I;W��:A�~60z@91���׻g���逥�ւ3���d2Po��p;��+G�(?�l
'7j���=��RR�H�G�j�Ӳ7h��N���6$I �%|���P�L�}��!��1�}�[�Hga�#�Ơ���7���zs���7 㵎���\L�aQ|�-\@U@����F�l&L�����xi����5���� ��>a�J�̬�0���$� ��v��T�����r�d����P��`�R�|3*U����t�A�-��g�>6�VAa;�P/�;!F��H.���'�ܣ/#{����hgZM�p�p3H�:�4hd��2b��l�KL�'��f.�v(K̉��
�����ݙS�.K��� V�v��|��1y{��mɦ�k�>S�����B��$���*���
'�i�%c�?�=&w�u+e�v�v|Wك���,j�䰠�j_��7��r���^	8���̔J�ǈu.U��`���{��X��'�`|?����tr
�:�Yy᠙�K`�!>z.��'�����]�L�?G�d���j���J*>
�nB�j������*.�m���v�:�C��6� �?#��	��1R��< ��M��>��ӌ��T[�Z�lQ�XM��uz���۫�5&,l� yo�mQ]a%�@�ґ͈s[D�+��;�:���Ǚ5��^�~�n�/�e��|Z���(g5��� ��Kx083�캊����(,B�bM�c��|*�L����OnVʄw��4�Jo�:�17��۳{��:���F)����=0�fP�/�& H#=%��j�\v���v�_΅����y#zh<\d���s%�w�
�¦�nJ�Ʈ:Q;�#L����-�8"cL�V��2�H������!ӆ�u�����;F{�E~�N�V1yw�dX��:���}jb�q{��0@�n��
83�a�i���>z���rx�JHx⸃g�]�����*�.����,�vaK�V:�J�c�������� he>��b��;�A_Y֪�:qU1��b���{�Bqvh�]~l#�A�sӪY�B#��(O�����4K��j�-��B2�,&���+Q�C�u��ѤݷzNq^&Iؾ��/.-��~o1w���5آ��� Y4�/�k�6p�r���	�
���N�*m�v)A��DQ�r!W�ao�P�짢��*�'�?�y������&��SE.ϝ�9�M���dY�,����is���P�W��$ ���#�3e��Λ��{��2��v�����#�V6���G22�����?nx���x��X���.���Q�W6Y3.���nC�8Q��+�ͦ�ǷŨ�~���)��������8��!���
;���iGdY�:ǅ��(P�-wS~�s�>3�zm�s	�"٩��#�����Z�`8Ǽ�4},�"���*�̨)@.p���j;oJ�%P�q?��|�GH�^"�{��O�X3��G�?���z��X��9|�=KIK�p�f����Bt���A	]�w�N�4M]>t���=�����||�v�:jtwv���z��ڪ/Ѯ���l��Oye����{��ZdG���Y��d�j`f"�4�|*S�����=��c63W0��c?�U�,�d�;�m�Aw�0G2P��}uZ)ë�[��7�.Ndg�aK�A�zL0{��Z
�d�f��GQ��1p��i$9�O�:*�k�A�R{�+ъ���kC������b��2���w�mp�=@Ev���J����/�G�A�Vܛ������WiV]$�K�ۮ�}L3	�I�a26��z#s��3nfj�L�L�X� )P¼r��J��~~��~���T`^��)�UЙ�ľ���Y+���8�P"e�e�d3䊹���L�n(尚S!��p/�A2�{���?5�Q�=!%��
�sK�A�q�>�ͅ�s��)���1��z*gX^�_8�C8���IDΡRy� ����".�	�B����]w�v�Բ.�/���g��	:���]�zV�R&���z���i+�#���e$	��(9K g����.��$���x���Rv�q )�CʻAnG������� ,���/�KUȩzVW���7���Y�y��O�T�d�m�;S���L�9o�F���4�U��&e'QI �*�h.�!�x��k���,�9��׿�(tp�r�(��
0�b�
�±`�z���AK�:���1�G;���KlW+�zxՅ$��`>)�b,7%}}����9+%r e�c������*T���#�8i�R�ݭ(]�y���lՃk꺰C��KR�9�;az�Vg��洗��-�a�I[�
09s�Iq���\ A�žpXwۜ*�.���T�"�b[L3|c4�v��`ζ�Q�G�G�N�.�%BB�iV�U/{�\B	�l����s��E�Mx�k�(��r��\K���;)ԞMy��Ո�K���fm��·�t^��}t��>
]N�ga�A0e0_젃'4�탣����zG�/2��<`!�7�]��ٙ��g�gu�1T��kf����ղe!�(�|����nLCe�V�@{厴���c�a��5�|�i{i��u���-"��,Yۥ,�B� ���ֹ��>�/v�5GWSC�fgPX�M�?���y���g�Q�A�ƃs�@���P��Qln;��0��z�"�c�o9�/��[.=9�����T��j�YŻ��Dx熘j����G�l���@}�-�Lu�4\Ypb7]V�S�}M!:V�ZRa�QZ!X�I��_ۜ?� g��[�e���8�{ql&Y��8h��p��
Vf�p��+��j�L2�ߐ%u@ڈ΀����X��nѵ�/ٸ%&�_S�g�	o��ak�:��/����fm�u���R�3�`����$��~(5a\���+r��#F���7qE7|7�*#��g d��I�:��G��oд�<�l�n�L�&|�o�%X�Riqw\ȬC��\u�G�Z3-��DH3.$*�O�:e�WT|��lͽ��	<���:�FI;z��Rޙ���s!�!QL|�o����P2F@���-8���d�K��w?�^��?����y|-���#9e�s��3�drLA�A0�<k��a��}��
�ԥ�]��b���z���=N�W��`�H���N�*����\��|!^	2�4wz>D+�M=��M�b�s�o?��C.�����Z�EBK�3W��n�odȄ��T��1)�)���ʧ���ܻ�7rK�D^�_qF�q�վ����=� ��e��vX2e���K�:�OX?0BB�+۱ص���ru�\�@��P8�X�u߹��d����m���
y���&8wM-�~t*�A�sc'�o"(yH�������}�"-��j玆+�8��7WH���(y�.G���U�� *�43�O�N�	���b*G����?�=�{�;<�!��/�d�b�!W��������rF���h�� \qq8ƾ:f}F��}�L�� �]9�R\kW��ubmd?l
��@��6�¾O��r�X�ܲ��V-�u����o��p�"|-�0��S5]�$�hA{rME%>��H��[ BɅ�-���f0�M�]ޭ��jRƚ]g��g��[%r-cH���p�D�X�3���&6&M�w���Б�]����H 8}AD�Ն��9�z��.�؝�4�1<%�O��c��;F+Z�{2���&9ۛ�
�yt�żȠz�(�3S��"�j�2Z(IT�dt���|g��H���4�-���o�J�<�
�Ťd(�H�E�(���s\e�97�Da�+������)뇜i�tHQ?P��M��g�~�H�o���*wiR� ��ϫ�ьlޘ��{u;����q������Q�&��S���[����Ï�k���2P�NyH@O�xߐ.�H�ik�lv�z�YJd��j���f���O�Q�g�aû��c���L�[����`�	8���*T�`��d�����XєGw���kG|��������|�L���v�%N��a��<e�o�`���a�Q�Ϣ���F�54����
�עp�T�G)$P������x�/*��

�;;�h������N� �N�)�6P�3܃����|:�Ha��M*�P����9�Iǌ����xB�d�c���w�oN��R2�*I3]�N*�21u����Y)��A�R�����w��R�0���"����r� #�,P?f/�nf�t˔|۶ݤu��D�&���D�$�zO��ŋҲ���8�U�f��p"��&' �x��߅�uKeP��y����
����� �����6%2�1�cE�}�9�.���e9��z2�ϫ����˃O��B54�
ᢅ�;ϱ���x��!Zm�=�ԑ%@0���s����P��k����#v�LY�����h�l�h���/1ր��J@�|k��C�aLؠp��x���o��Ui	�u#�m:��@�~�h;��Gu]��!��-9î�r�Ѷ��C�?Ph����˺;�2+ �b�/-Ao�v|e�<L��U�#Zi�eE� ����h��V� {�U�I�t.5��h�����.�	W��E�,��кs��֎����6��}T�q	=#����!jN��M^�ֽ�̓��w�\uSnWӓն�;s������J���,�������齓�ra�60���V5آE67dA��� �dJTɎb��!��f�h�,|�)����LQϨ�w�0{K����/��� 3o���9
mxR��}��#���ۋ<o�zڜo�ȓl�Vi5t�Qo[ڤ�F��qW�~�/�hs�^��� [].Ju���d$�%��|�&,��u7j����O{5g���50���)5���eq��F���c�>-BDG�e�{TW�y��TX��3ʿ1|�S[�cJ���e×�=��he���xU\��G�M�:+��3FY�Nq>��q�7�d�iB�WE1��U���g�Wm���*�a��+Vky����X�Y�h��a�#4���]V�@�2���eN?�8�i+*OE�2��c{�+XP&G�E>�n�3�i.Ķ�	�Q/�g*�Wf����|���3��T;�kO:�����>�}
Y}fd�[Q�&y9��8�o΂�UH(_��*�vD�[��&��xA���^w���]7t�z�J@y��D.+���y��h�����W�H���Z�CI3�S���4�m�(L�z�tb���a���0z;+K�R���#Bݫ���w)P���:��zJ�}
��b:�:�SA���Tr)����\����դ���b�H���T u�3������������+�<S�Zr�3�����]B4�M�cr �
����>�%y8+��c�Hz*<�������ab�mr�DV�
�4S�a�'��'��Yf�gBf��N�����~%��2�	S�<'8�����E���g��]��|ذ�J̺Ti7��fئ�Bm|b�0�C���玕�#�r��_��-D���d%_�o�E->�'��!&zkocSx�����Wޥ�7�h`A��[7\�1�od�̮:X������e�S T@�~���N;�#��&������/�#��}���Z�P�#ɋi�a�=h<���Vr��!���C�O�/�����y,�J_Ad����1ú^��o��O9��3�o��醏�a��#�ed��Պ�_��*��)�^�g�J'iYS���~�t��*C��v��$+���t�ji�(jIM�h�"\p]|?�֯N���#�]�!{�?��ϵ�Қ�J��G@��8��������h�c��l��	8s�S�V'Ee4`N���|R.�,(��\|��}hBӋ*��jgL��4�Ε�G�0XP#x*2��}o{,0|CN6�#ݫ����>�ǹZlᖘ�K!X�8�ڀ'���A"B�k0�����i�Z��ق:֝;�*�Ʃ?v�_y�W�}^�4���y�1UGpnz���@>(c��32��<��_�:!��˾�84�D�4L���߃A�ĠvIڣ��>fh�~�q��6��j�5�һ�Ya�0.�s|��Oթf;d�]��J����I�]�.������~9��xąm�����kh̟��!�˯�FW�5�eov�[<�s��k>���2wTa�1�șBm*�5�F,�,�e�t�38wuRgaOS�֝b�g��`o�7�βB�����߅���u=[�%��JK�7Iø	��]Jxfh�̞.��	�I��`Z�s���=�'�pדy��c���9J�Q��T�:>5���{>S�Xd�F?��-��˫���Is�&U^hK%�A̐�qm�=���`�X����9�/g?�dୠ%����q�^��%b�-.Z4���^8���:�҂'fk~����C����x��ա�l�R��s��;�Ju�o���&xw�P=%�NI�$�TN,�q]��J)�� �菗t�L&0:K��8SjS6�|i[Fp↦q�<*�$��	q|K)�Rܟ�OO�S���ms+>��ky?o*�;_��8�*$JX��vǶ���k��R����jX�db����>�.��ook�L�-����˘�#M;mFT�vt�cU��Լ*Ǥ�f}V�D#O����fm�#uEC�W�D���j1�e�*�㛵zkd�ʡe�����j\^��=��q�61��/����P�ݼ�@ӌI����!i����~��sk��%?��%��F�&DZ�̅�R��ǘ�WbXc�>T�י�N���)�s�0�p
8��Ђ�20�1�@�H���Wl�daߝs�S9�щ��|������S#s@�{VY4�f�©/G���?��< �]$�uqwE���/�C��>+)�ΕI��><�:C��T!��+o�H����c%��6A��CĊ��h���2��x�9��.�A(o���2V�}g�, �n�V���`���2ͧ���vBԵ��m7�́!V��?���i&����ʔ�]���ڙ�=�p�k�]Z���i�[��w��6�h�k{���:Mt�H����b-�C���fu@iLv ���Á)��B�����p.Y\M?ן�R"		x�-G�m;�f�$ys�V+��5�����{q�����l�m�I��TlX�N�����ZY�݌;�g\�/~�8[�0V޺�^F�rD��/��������9p���nԎ}H@i�}�*�" }��d�~�i�����4��1��Ñ�6ӆ�Z����X��i�G��lRӥ���1��i�Q����3���>���xBR�s�Oޯk��j1z�$%v	�ń.��"���E-hx��K��&X��nP�d�=R8E�At�n�䏉��dR�k���X�ﾛ�jv����_�:�0"�0�MU�;O�@Zב���mB&��T곂�����Q|7(����@�Q!~���6�S`}}��f��Y�)�|Jn���[	(����M�Yqn����\��٢#���0�<��:�����F��X�����R%P�e"<�X��w�����=/7v4�{5Sr����Ѣ�H�]:Vﴎ��
�c��3
�P�6�d^6vΊ_�o�x�b��_����5�W-�!_xq��tor=�i&y7�rS$�Xf#�����gF�D������z��ZԷ�J�OD��{e�
��x��0pDio_�Qe�oH&���n`�w/��Q�~�p������+���4y������7f�0��Չ�X(:��Y�a�m�q��U���N3��А|žHr.xa��
��g�C����B��&#�h�ТU�q�G�FKc��'k]j�&�;R�ilS�ĊW���ݚP�^:�+u�󼌑Xr�H ���*�.���h�,ͨ�T�0mc�1M5��r[�I5X�9lu��c�����g���ED	���ԧ��#0Z�"ܵCJ��
���.g��[��-#l�׉_%�vG97V|H������[�j�x4�������~�`o�k�W1��Da��&L��,4'���OQэ�#�9Ȭּ�
Xp~VjE����8�R �#���Y����r0�mu��^�6Q�S��@W��a���O#��Ef.ԘO���_a� vd}!�r�����+���� �B��P�[���WL�
TE��l�[/�>Kc
ã���{gj���,�MaTy^+���+4i���C����zu�&K�Ի�X�)2�[�u{��&t3�Ü{Bwoӣ����+@˩*�'�;���C�����&o��KƑ{�tՏOܙJ�rG�3}/�����0�w��pG=4�fl�X$��F.kԮkBg��!޽������4���ߟv��s��Gʧ�6�bz}��:��ZR
����X�buǤ.�Xt�{J�)�.�!�C@M���O��zc�'�;��{h�19u*��a�d�����C�g�r}琑s%�~sKEᵌ�������n�?���B47�.7�C�&\k��n>����}"��f�\�3^H2�C�[�� �gC��͸���L�P=�Q��#|V3���S�z�[x�j���k��k�ʉ�-�Nڞc]��\Lء��3@m!c����WM�(��4�pw?CF7Y��)
���+v��=n�Kq� ����0ms���JA��FSW�I'$XL�1���s�B{۸�Y����E����5��ă ���\��?SI<�`�^�!�h�)����Ĵbiޕ�#k̵�6a��z��i��R�t��O@t29�0Fk�ܽ�f�1���o9%�苊�دp�q�d3�([]n�c9�2������R��u�'!hƋ���vhgT�`U��Ҷ��._am�q��8���au�ٝ���B�ޟH��q�'�漊�*lv(�(��"�3�Hp�ۛ�β �M&-��=�^
p�Ep�<��t���P_
�Bv\��Z��?�2sƯ�d�9wj�1��/E�\G��! ��2Y��oT�����=�=���.�BJ���/Ԧ��0@	~4-~�7�� �T�㩩'��Lւ���>�e�A'�$������A�ܣ�Lvi�#k��LIş�x/��de���B�%,��^��4j�¥� |V&�<����x��q��3�<`��V�(O�u���@��Z��9�#����)<>�蝢@�%�>k�C���]��]fݝYg�_L��[��-[����;r������u�����c2G��⊞�A�Ʊ�G��]In����\�'y����xzCze�%" ���l$�"�(�[R����/7B�v���cE�ۥ���|�3	"�wT�n2rۿ���$d���:�<N������j�w����g��8=(os��G���A5o��&�=F���ٖ�e�0X;���ey��̴<�Ӽ�PKf�%�����6�QZ��������`���P�_�Q��bYXu|}�,�a��m��{CTJ����N4����jQ"Aw��o��B=[ҟ �V�.�M߮8r�O dMu%�|���Z�L���*��	0�#7�N�!���ZԵ�V�'��"<���o�q:ު���T�����	���rTI�]%�r�oU�ex�K�5�,y<?��a|����~)A.���ە�74�n~�.Ѯ�x�G��M: �+2�>Ϥ"�����_�N��-4;�:JJ�������>�_7�����h�Ò����� S�����jN&G�0�IqC#5K�u���v��h������&���>���A������ַV .�T)?#�3�ėȝ�/�<z[P���]�zjC,kd�YLm:�=�
z�}݄v^�7��O���`c�_4rxQ%����I0��c=�_>X�Y�-�.#^,�{xs-kY+���2Q�)3  �������K�F�/XF^8�EI��^^A��Q���˵tG��"�q��{ܢ�\U�.~r��1��ݦ��+��N���(���S��������4{uQ��P�;✒h�a�B�CCݣOnU�zr��n�!Hj�������\��6����[�e��wLM�w�<M[�'Z�{{J����ߥ@����#��X� _�U�z8pPIj}EE\�f�<�<Tyw�0�8�d��	�i���j�?���Qkw?�V#��Ү��`k�7m��hM�(�*��\�ܔ��u��aY������Ք]u�
;p ����&S�zs$U�G;�z�W�H�@W��<0���ԥo��kmC����ן��ځ ��c�>Ew���Ղu�r����2�@S�� �Q����n;|8�����k�D�f_/�HT�BK"|�l
������"�)	�jH)p�z���T�M�h����3���,o]&�%so�3�.%�0�0��fOdԷ�?�J2l�J��KYlh�J�Q� �=�n�]�8@����N�T��J���j���{��������>xW����S��M�Wl�F�2qF�QG怖o��=���(>�Ӿ{��w�$����:T��@a����c��g8e����tB��N����cOz�5�t4'��dS�{�yP��~�lMo�cS���H�ç^�w�ż"�|�%� =��U��eE�㓐D2ץ�t��|��L�GB��od�������,�*�7�H�@A����uǤ%mn�7s%ύ#��>d���"�8��j�3�$� ��,�4B�O��٬�C�����g�ʆR�=ZE��2:�?^
������E`�{M��M�Wő��.��l�TO]����Aw=�k�SW����򥌢8�Z��,�n�7���Cw`��_��ʻ�-l����)Ҷ���e+�r�}e�(0�1�����&Wj�r����`��Rm,<j�Vӈ�G�waG�<e?6f_���Ҥ��!b�D�0�2,��ŒnG�%�F��&�`���(I�M���&��W�6j���vx�FU:�9�3��y�P�_�[XseB�xA�0Լ[��F<kj�G�_��e��W�R1]X\�%�7ezG���WĽ���8CgT%
�z9�b�n����:������~A5��l
g��������Ef�U�X�f��e�05�#og[�P�NZ��jf?D��lPe+Q�-�$4Xo"��\x�H��B.�P��ޫDޡ����(ᑇzq`H�C}����(Z���*
Sn,p!�4��I��5O�`�P��O�]�z��
M�k7P����L\�2w9p���i8s¼������!��p�Yy$�/�$;ϑ��K��Xj�]���%����t}�L�;@�����7�1�s놋I4�5���0���=��T���Q$QF24��]��,f����aUлع�@w��p���j0!�jLD�z����ҍ�Z:F��A�Gvb���[�'7��̙@n6�v^�jZ���^?����,1�^��׍��*@������m3�k�1㒜���r�@�z+��*�2�$���bb��TP���** B�9�a���L	Mz� *�δ�C��QU!���'^uy�T�af��R�}.8��X�U0���Oy��ڐ]۫n+�t�6���}���*��3����g9�޲��w�7
4YI-��7zwȂd����P+�Ἆ<�S�Zu�1�ˏ#�p8}�eJ�E�����T�!�ڥΓp �"��I$��? �7L�[��~���\�?�oKtO`��r�Ā��4.�S@�@+?*�;`ઃ�l�Y7߽*�z�N �j�F;-��ܢ����uꋗ}6�P$���Zƾ�!z�?�il�+��WRq�f�Ǭ/S�K���k-��49��]�N�^ԫʾ*%��������{��&�%�pA�uZ���rk������*L�m4��x�'���6����{�<m>rF@���8B[ = ���!Q�}y	���CṊ��Z�fr�FIXEcu��&��:e?�Z��+��4�H��S^/��y�$
bPq��Ў���L�^OЬ<��Ά%��d�d;o3�����1ڋG>��T�ʉpzh~$��S��Y�St=�̟�}�:�I�B�����$�U�z��h�M;`L�ѽ��]���[�ä��Ž���PX8��G�̬��Mb\OѫB�2<TPD��ӗQ0��6Y�(�W,�	t�_��]���2��yf��:��G�A���ܖ�
�ez9��
A�{��T¿&	'���{�]�~ş�_�e�-�z�5LA��NvpU���G��l�1�cvO�<�yH^;|PnI���_�z�S�txAe��Qn,X@$kRςg������^HCrI-镹S�-����D]ya�K=
 VKA��Nw����.��tl>�4u��̱�`1on��;��i�G�r��0��^ӂ�"w��%s��Lr�<i��*�ȷ�lp{���@c�
4Ϋ36���jr�o�{�Zd��q	lD����=�4"���@M/�f\��=��8� Zm�#N�t�I����8;�?Ƚ�XK�f�2 �3vִG�lV�e�MP�A�~Һ}������J��1L�Ҋ�K4��*Q��l��;�����S��Z��R��Öoy�p���3)5Ȍ�𣅞�~��O�w_�kj��˦f�L�Yoҕ���s#�?m�Y�����V�*��������^��6�ZTE���<�%���J���������L�v萙ESn���h��C�K��f�E0-S-^���j�T���=z��\��,i�]�}�uH�Iy�_*�w�3��c$��B$�&Z.�͌�a�S�
uN��M2�Ğ�5�� ,�HeE�	� ���`��H�S4�0��|���Kk�l��s�`�0��S ������Ff��Fb7*E.�a7|;2I���m ��.�h}�P���ڸ�P�t�LT<8�n�|�	���X(����;�#J����\�5�����0-N.+ѥ�뼅�dy���Tɹ<����b��a{�ƢY��O|����Ʊ�ʨ��}�d�U��ԥ^R��X���b�P�g%B�C����2��zO�x����*�9��u�&*n꼵��_�ih\��Y�؀䏎J}j�M���Wy�݊��c��)�O��y�?�O�Q�Q�U�y���/\�6]s4�!ʬUv��-�m3Zrԩߧ�*���[f3|-�筟�>�����-GL7��@<�1p8���f���	i�+GK��c����j�vd��w�ux���NC5�_H���j~�R�x��ݹ���ʌb��x������C�Eo!��Q��
�¤���p�w3�K]|ܢ ((d�s.6�>3�/&��Se�}���i��F:�6���3��a4$�I#����������'>��D+��BZ1+���-��4�z���-#���n�Wh�`r��$��	�9I�1���AD��4����2?~���e�p�(�'Q��ȗR�|�A�n��T�Y���נ"�~�m��fƨ4$wԆs�s�MWd����U��1!��>w����g$�^����'on����D��mQ(6��_(�k��/+#���j���(,WZ�^�/����1����ߩ�?-KB��q�ap�P�ＹDnQ�Y܆k��؈�=
��K�#��Q��擄���� /�Vm�i�����.y.�T��m�!� ��)Np��Ӊw�]����G.͝���VNdGd�b���� ��ڞ�˝�tN��k�KɞB*Hh'	zJ�3��%�aR�e��+6н9��D}�
����Yu˸55}%N;��I�3k �?|v��@8�
��#�k�0V��Pl��� �8;$g=��@�ٻ��M�:�������=5껷�W�^7�l.Ң�M�T
sj�i  �nya�X��$����鎾��8���|�߾�F{�d
&���iO�ħ*!+_\�F��3�{�߲��.�M
�X��"���)&�b�i���!����"���oH�|�Ψ�v�.�>��=q�Tr8�q�Y�.G��L���+xg��T:���9Y�E���]T�h�ɵr� �T���ܰ��/@oЊ�l��$idU$���Rӷ�%J/}�|j�q�\K����E(�T22N�"i{޹�
�Y���J�
����tl;g�r|%��ɰ�Xv�Vھ��T+]�^�y�R���.~jH��ٳW�"�w���?�Yf��<P��k���&�@u��U��6�'x:��DodZ�5a�1A����a
Ͱ�1�~�7�c����Ҳn�Z-ђg��^�QrG��o�8�ܽ����l2J>�P� O%��хO�M%��a靊$�݅vy����|�Nzf���|̎���y�_�t�M<�ave�@�ߓ�.�P���nZ;�
+|n�a�
?��"-਋Q���@�n3%��:��yt�>A���_��ᇈ�6Ӄ���b���h�	;�Dx��	�,� ��7Z�[kڵ�wt.�}_�YI.p�79��CL�"���@dY4ow��gVj�n��������[\ˌXZpM��f>FW8�ȱ���MZL�ph�:�7O%� �3�uGL�V#�	̵�x̞�cn��i������+�e0D��@]@�:��o�m�HNE�)�-�����l���������M"�ii�C�G�	�<�esz�[���R׆z���b���0�j�����{k��!7���f���D��-������M����>���������&�͗��U9{A��a״'�l��&T��y�����Yo�z����(y��	PN���(���[+J������bsf+Rr�Yc"�2��d�@�����:�"�Tk�(��l���y	Uv�,PX�З�C ��SfA����Ǽ�f*�N_�*AV�4B?6�wٺ�i�x�ȷz$ ������l��DD��ʏ����hq���6����5C�sU�,S�/k�vAt���H-;7��b���O��m�>�+/������e��iT�+������c�]�!z�����Ч��F�a�7	�ћ�F,˧�����E��܄�9c
������iJ_)E����&)G/��C΁��|��3�p���<=�dI-����ك����T������!�w��P|uiZ�Z��ؼ�8Ӌy��������	��J<��ɷ�zi�Ɛ���'��F�#DP�F��9�XY��&��3��\Š�R� ��3]��i��ѩ5M=׀��To�>����i�s1~*q�1�_��}~��9����&���q�j��Pd�C�y0�cً�b]|
a)�$�Q�u#= ��#�0h7�D��u��kb�s�(���ɭ�f*R�QC�3��U$������h��#I����V[��6KH�2&�y��u��
���{���N�ѵ��]�
�����X�����9��z��R�gg�B�s`AKk��h���M�\�lLh�(��d}}����r=���w���������s���.�j��<��:��,��S�"�{�Ⱦf��	�'b��C��pzj9!g��Щ�z��g�do�|�v�`�������S�����K�b�q�+qU����?e��@�p��rT��Jä�4ˮg|?��W^�"*[~�=��2?���b���磆dv�I5o�zN��F���x�f� �"8��3�a̔t:sT��EsQ��&���Z�;D1�W�)�2��;�k�4��p�Ʉ-�N�����nm�e�V�9w���w.�ԩ���A�����??�5k����(��Ko��w�Y"��+u�q�g���}�Q�WbD(����_^_��¨���A�c��q[1��3;��h���ɰ��?Ĝ���J��dA��Ҫ��@[a)�q��<kK���z8�X�c�l�=����i@�ˎ�h���0>���--����˼1pDkR��R�"T�sZJ��9}�В��@�����.�^���s����v.�?�nT"�>��r��yE�3�Z��i����#O8�lbz#�W��3f�#�Nr��9 % �?F��V!��}�Mb�9�3=6�g�H��˵���qo�DA^�%O�I�Ѕ��zh�x�3�R?����H����,�4�_�7z�H�WX�ڷZm�kJ�}�ǆ��*,d�u��n�Գ�~?.��]�����/�����[as��q� ����i���S��Iٳ�1m+�X�x��̠N���6j|����3��?�d�fz����*�\"��#A���Q�D��d�ݘ���}P��@?Xb�O��ZǲH}d����b�T�
aU�Ԙ���Df���ķ>$�rм���L8�SI&�����yښ��k:M�%��8�ȍXƴBHl'����c��Pu�`$���+�R�%���i7�p��A K\Xй�1u���{W�T)��\n`l�J伮?~Hk]c�q[l_�TT$H��Ç� ���=ܼSMս�������X��yV�?dI���(�mY��S<W���+��^;V���b���ɭΕϥ��O��&}��0�:�4�L d� 7$s��Xϋ�{c��D�_���r�׻w=)IF�#o|��L`�f&F���u�>d�"��~"���h9Q����[Zވ���a9�4R�	xDd���~���J�����$D�V�y��!0�SF/_�	�-H�&ꅔ�ު������g�L͊D����~�p�=a��{�_10wI5Xn9�t���ƶǑ�P�0k?�x��63�sɘ �vN�Ҭ�U�r����3Up!"�2�m�CF��z�G<}0X3��&3�G�y'b�v�܀��L{b������Y�:�S�V����O�3�<-��Yư�Tb|���?M�-4�k�*�-�2zg���e�B�?���~���7�`E��دCn�m@�j�i�qk]���/����PQ�����I�����M�:�R�Q�3 �c(�&���,}>���a6��Ҿ0�ƀ�;Ht�ZO���Q�~����k�=��
	ʲ��� D�!�g����5���")v�� G%�#����|�gķ#A	�Gc4ٳy�	l�T���t�9؊�!��A�B�����y9�����>��ψ2��t.����!�D���|:1�8F U��HYx�{�Ԋp3�A4�r�ń�@b�4��9TK�-�bؕ�������@'�ø���"D�7���ꨪ�D+���ߛ%���""R&�eJ1M�a�'�h7�da�t���@5�����a�]��Ě���[�%'>m����$��P%3�*� �+k^a;�y7�)����R��Ue�¼ӚE�Lϵ$?gWx��褎䃵wyh�JV�1�g��R`�7>L���\\^����9��K��z�D����@����s������9㡓:�W ����(-��/�_È�����eX���r���.8���/�Y�BC�qm��e=w}�9��wW�^�Me�L/A>j�N��-1���N%o�ՍC�h;�w�(���}ϼ#:��D�5;�pͻ�؀�3���ol��l�a���
�A��N�Z�l�Dܬ��;�i#| ���6tcˀ�������s~�jY7͙�{���
,�霻������'Ak$X�r�z���F��f��TX8h ~]�=:��� �����$�ԥ+-
���Q���5N���wU5���H^F���X���o5,6]�&IAXi�&X�j��H�<RBQr���5�9�C��?�S�"uT�سYVѮ���rXڞ�-���u �v������/e#-��a��҂Z4Uc�]آ��~G�`k�W-�x�1M>��'K��T��(�R*��d~�$��hL6뾍���ƽh��ǫ����(���B#YD;;���x5"i'�W+��£�"��|�@�vA�I�*DEt�_B
�\���Dz	����-���ץ�����MG��8�ܢ�5M�8��9����fB�fKS��|S�R�W��p�m�:-����@'PCq;kBB��}th���f�\|�������!��\xk�1�c�
�������#�nn��4[���� ��=���{�Pk�[֘�瀎�WV�Ǘi�u��^H-L�]f�[�r㗱t�/��Y[y�#����ƞZ{�%*3Kt��Nَ%a�FrZ `��t�T��Ė�/���L>���$3
������I�'k�%
� �4N���!U���P�
~���-�B��k��
�x�+��l�]w%������@�?����{C���O�ф���� Q��1�UC�S����:�<<��ΐa��g����3q+�������d����OΓWkm�g=�<O�	���f��P�FZ-�̣U�0��-��qF�$���O��'یW�I�R�\4�\����,;���u[u�¢d8ہ���v�#τ��Yp~��ѧ,�3�^+§�)�;�!n+[8j�4�0�%��W�[>�y�l*��1U�d>���-�5UR3��De\�v�a�v/I�4N��ۤ�m�h%��$H1D]�S����)N�@i\�䞓y��>Ƙ,[2��4o��x4��>?�W�ep��߃�9����6]$6�]tH��Y�덭^ơ#8-�83��'�Nل���*��Z�*ծ�R��A�7�����+�y��V^wධ���f.�Aغ���	S0��b+2M�pW	��.��)�:q��i�����5�����)] �	k͖ꖍ[�o�V��ؖ3p��id��k�
ԡ˗f��y�JtrǸ#��v�5���Z�����ưh��@��cώ�:��+�9��y߬J�f�Q���z�Wt�L�	��S�l��Ҿ�G��B����L��i#���?�URi�07���EΞh�}�83��AU��5<�玲�"�"�
w�ˬ�(���*K�6	�Jp��&w���'���v__e����ؒ^x����>=e~��t�d4[?��&���!F$r�c�HKt�;�o�'��ǣ��tX����Nc����"Q"�k�Ò���[![Ъ1����b�	0)AV��f�ZL�I��G��A��N��5�s�:H����B�f��}�1�l�H@��mʎ|oȘE9�C
�g�z%�M�v)֥����BQ��4C�S���/eePq��5�y²#�{+V�L�����(YB_���Hb�$b�Q��(���=J�␶/F0bN�*`�B<��$iH���S$�Rf�o7i2�}p����s�@����VF���M^׻����h3GӶ�R�SY����g
���!-�ǉ�ܿz���]����ɟ��(n�]%�Å�Ӕ�s���`�*,�&2i7狅�B+�z�����<�`��@C��VpH3d���� ����+4�\
�?:�x����?�1�*�,�s9yyM<���W�L�br���8(��|�_g���B��+�=BR�I����U$��5C����ɖG��g�s`b�gS�S�A���y@+%@���̲.Exg�b�prd�s���/���R�
$�L�`<娼�aea��I�ze�jv(�nc1� �p��R㰌G��+��O���វ!Kv�~���i�EU�$y����������p�vMԎ79\��d��2��^4�8�l�WX��zvŌ+CkH��Z��'ɐ���*���G��ͨ4�O���
u�ԩ(�/(�Uvy��Xu���I]�ԑ��" �pY:��Ҹ{{�V����&�#F��x+�Q�i#�>�T��`�Ү�-�B��P0���LJ�7'�/O2�с�G���f�ގ,�/97�ʡ;��vF����
w��WB(�X�Ŭ,f�%�n�'q��0���o�L	��f�d���7��근����J	�p�Io  ;2a��l���@�a��@�j�7���)Ö�w��q���tr?miyU	y��N�L͖���P��吺�ǲ�Xb�������B1��m�E�S���a�v��`�5JV2���yF���%#B;L�)��W:�O����r~��z�(�>R;P�{�Z2Cqo����0;��a�t�0�F�Br�N�hfzI-�۠�8ԪJcz鹏��u��C�C1ntC��\.������_��A}&'�O��t�j��=z$:8V�F�㣥)���]�3ߴ� ��_s=xJ}��9�B���)���_o�s�����-, ;+��
y��Q����[C�	�5 n+j��O�졃�8tw����+�tdS� �nЅ�	;٫��du�(IE�S�O���Ƿ��|&��}�<qf�&����\��1e�'N8�����Eӡ#�1�B�Ȳ�4;�p�}7�����(pR;~�F~��f������KYN�������7�E���W����&�4"xM��W`(@�����DE���wpk��O�<�oº�*�w1�@T��b|ї�('}�{���a3d�"
6�O<X ���rW��%�����\w���E�]Z5�W�l�H����G31þ�V�[�gl�O�u�
��D\'�����ފ�'s��l�}�8��R@Щ�x�[�DC�������1X�8 Q1���mR��VEĆ�}�:*2%�l�.�}��I8�6^�T�p���Z1FOz/7�b=�m��uGk�W��WR�rg����u��r����(�#R�7}�{G��$IA
�@����W"���M�\���6����݃���=�w���|:�Z���>Ƿ=�Li�1������<s��3m��+-=�n�0�n�Ѩ��ܢύ�H�h�ghdG�?����?^��:O|͐�e:?c�ٿqΨ�k�1��c�짧?��5�q}Y�Qo�Y�P���c�qV����,��N_v̈n�y����Ox$�5�d�V��}�G�jj/b����m�RW�Gb�\pV�z��܌�1OP�����V���O��Tov���k��D�I�[G�4�5�X��~_=�r���z�+�ҩ2Gg��;}�`Lz
Ӻk0��3��\ּ�k�_�*�G߈���g�D�j_W:Ik�jb���G	�.�OL,�)�=������r��B/a�vx����h�tX1���.���u�Q��7]V�4�9dR謦�b�,���Oߏ� ��Qe�S�8o&щ�w���U��C[�$X9g�毡ӏ�^ ���9�����tNr�ېX#�'=��^���6�%�6�mPG��^��S.��I�^{b-'y�6䌈a嵽vz~F��{����� m��2��l�z�P]�/[E�Ke�^�Z�	yWh7S�Ͼb�yt�[�Z��,粆�O��G��-��&u�� {���~�p��%E�SY�$��w@�(B�}����gy�O3C#�{ǧ�C[����B�i���/G3��]^�*��ZS�^8���1�Al�(G�v��
B� �<�)Ik�� ��>Z��>N1\����� ��Z,t[xl��S*8�b�f�SR�����j�'�0�k����f�j ��5�r�)X����nMt�Y{�M�sxR^�u �u��A?8hj$��k_�r73 0H\<P��el�c��٫�[!y�D�L{�Z��	ٓ�K�o=��0�N�-'���>�����0�ۿG9�/�w+��r��mj��m@��/� � 0q���`^P��,��fP���d��v�/��Y&i� ��E<sO�~�y
�o��QqV׏W�#\��1�P�����ZgNJ9u��4'uP�KqG� �b�2u�Dٕ�#�`�7���⌶�!�7�,�:*W�������K�3��[�nx_VrZ��ӛ�/���V�:�r�R��}�U��XXr*]-���)~�c�AjDd��R�, Z�~�4����[��^�T�Kd�N�d�ӝ ��^4����E�G:~�n�Э2ظNy�'��߉,���7��lP{���sQ�|N����!�ډ�|�$��h!�5��C���s�T��&�?*iV��/����Yw����������&J!@b�3���v��x�SQp*�>�ܛ��0Ma���y�i�Z�mը3��w�g<<�$s���]p:���" S�l1GW�d{ր�Q7l`�|�+�J��a2ݻ��*�mg'�!o:J�_ r{s^$6ݎ�?��έ�Q��9���cD4߹<#�^���-(Ц5�<���S���HU�J<��ޠ6;,݀(��y[s�G�l��%��-y�6��ؙr�dy���)`�\j�N"�M�6%$K�>ޟ��J�t�<��J43z!g.�iH�̟�U��=E�0�Ԋ*���^�U�ɩn�ዣ����,�e
�NL��sM�m���0����,0D����2c�%��H(�����F""��K�:�.�B��V|����7�冡d��:��K BE�T`�03��@�c�?����e��a�֧{�4N!�z�+y�`=Zs����*ˮ􍺥�}7[�A��{����������)=�K�L��S��R2|#
�������ٙ"���a�X��/y�,��� FW�6���'���Y�i�-�C�:U���4F6����=)貮�,�����1��^*jf~��' �P�`W��h~P��8hK����5�}����e�ٟ Z���>�bA�X����R�'�Ij��Y���Fr�Sh+ 
�Zl��N��b!�of2&���}.�'��N>.�?{��ɶ��D�#�0�������bH�K���G�U$L|~��p	oҀ��~���S�ץ���F�����l[�9	'�#M��L��tŲ뇘�-��>�� tAz�O���!ZD����+�?ˎc�"����F�Wr��NCM�Oj3W~�8�}�0E쯬���Ie�U�M�1��^���R��xi�:�<�6X<�v�t1�;7�Ţ:T|՟}���\^�b��5fYgmw���4��ȗ���������x&
X97UqSG�0�aR0O�
����첓nC�<Hkހr�_��q'"���P���Yd�5KTV���57�1��x\�Ӏ���Ф^��'�^�x�I���n�]�1�:~#�J0 �8��5r{!��#�1����ϻ51a0��S���ջ�e�~-˃/��O�-!��˝���'L(�<���7z�A�މ�x��:�,R�Q��/��}�FM�Q�ԱM�[���{a?�qY���q59D �u��t�̺'�F:+�{�b��З�[�8��W�i[�G�Gq������=���ᮘt��-�PCiy`�+��&��>i�.���
�=������.��5�1��������c
�%�L���`��M�qm���d����ԣ���Y�֣t��jGbi�c���v��������Eq,;Z��F4�Lp	[�LĐ�ۜ����l��P}�i榈.�>:�]FՁ� 2����K�VJ��:G�ܦ6삝d.��!Ȏmsw�1����_z^���&�n. 5S,/E�I����<k��}��,�T�^@tT��vc*��˘4���~��'|�[g&/�t�����ԜWi�	���g`5#
_���&�ߧƥ��G�rh���t��#�a3'z�t�1�����$���+/9^���38ڝT!E{j��ܒ�ny��b!ǎY�g�������������~B�ቂZe$AB�v�$˞4�]�O�C���.�x��m��m֊��nt���&m�eO��{@`n^P�vL�)���n�L��d���*����j/*���>OF����RU[1?b���o�:���J����Cg��g.
�� Z���9"�����B�D��Ƴ9�EzE��o��".�Ց�5:�����r�I��C�7�J�����p�}�0^�%���3Іwr��[ �?�g��X8�:lҎ�����p!�}�Z���Y�)��悉DdV7ҶK�#�4��8Cn�"�,��JS��m>���켈~`=<�_�]�<���[ޔ��(�g�:܆�,׊h�Đ���	`��$��lz�I�Z��K��3�����,qm�I��s|�bH职��З`3��?M�%��#[5�B�R�ӀS^�O.O�<��LB��Q^�c��-e���C���O���kkrEIJ�sA�c׽E.O�|��\S�ϐP�;�J���l�A��C�_�N)�PwݽE�]�ڟ�̲�9�b�>��F�O�v�vb�.X)��{��K�XSJV]yí|�+�9?�O�(C~!�'�p�l�n��$�Z^i
���u/tI(IK6i�Ќ�_r����������]�y�@���H�럍$���h)��"�E�Y�\K.hQ��y�W�&�o$�,��ƚ ��1q��D��;L/G�(�p6�Q�fq0NlZ}Y��ɻ
��!oV�,7�o%��U�L�=ݹYbdJ�w�㝹`c��ۣ��E|�R�\�G��O��ix;o/J�ᷧ!r�����e/�ٴ���T��٧��;��+(�����8<�ur;,M�oo8��)l��%���%S�-�ΧN=���ؕ�]^�Rz&�?^O�x{���u/�`�@���������!&f��xrK��{�6�q��R�������M�?|W@��@)*�5��4��*n�U���P�13��5h[�AT�nI���^�����ʑ�nv�/b���L�
(�^�y�x~UV���w¦/�=�b�}�7��*���%��UȄP��Mg��@�w{h�s���b�����(���8��0ē��JK����8�_g�XiV�&*��4MC�S苧��TP��(=�]�jh
�Q�0!�Ӑ*���"����N!�?�+�� �N0-�'\-�}�R�n�[�i���h0�8?��a��<L��0U�oŤ�!��-��;V�z�1*��z���$��~}�c�و�Z�������ڢ���I���d&~�\`�lo!��K�̯��<�Q��X`�<i�'κj���27����l��m�G��R�-RIv	u�N�B\��9�����)z!~c-�1���D~��Fz�e$`�h��v�I��.byժ��:�����Q	�'v;ؼ�iMN%gC0L�d�2��j��a�X�5�R��	S�c�n�?�m������7͆X��գ�/���ەS-R�α��*Zt�U~�I�P���ô˅��d^n�����C������Z�b~Pz��ұgxJgG�$�J�࠴�_�.�aB֕�8�W��9D���Q�T�#ɜ�+~�a�P�ԁ��57��ΐ���W�_��h�G���Y�̳<󨏘B��[�S�=���QS�e��*kSyF���S�6�o�.b��'��:)c���f�ǐ�2�,zQ�U�IJ�e����G��?�;�KK�P��)��&AZ�Z�2x��ޘ��������C����p�"׹��$�,�'��ks{�=�x�-���|FP��yK�"����$I3]�/g1�U҂���Ǜ�#���=D�U,N���TuP��{S�E�4�.�f��!J/ſZl�[0-\=��q�I7!aGJ��u�F�n[ru$��[�IHh�&�y���f:�'s��4;���v@���Z�6g�>hA(����;w��j�eǃ�	�=���.��!���OZ�W,x��F��%�2��1C���BRƆ�hL�\�~_!��z�GS��~�����{޲s�t��5���Y߼"��]_��[�:�)�f�;��.�^�	ŭt(�{;�4읜0��T�b�a���Ծj`�ئE�q�o&���?�	��K|�J֭=���چ������ӕ����w�l��J��Nv�Ns�=eW#8���2W��uV_�QQ� .NmI"~�����콝�n2�a�����,�r�4�����ӣ|��#H`Bۘ��}^΀��B�vXh]m�� ���O���9��~3cH��u/�٪�O�����4�k�F�� �M�.���7����@l�.(��2���*��S_q�S[@�@³���Y�������d�n�Hv�A�(�)�f�J�.5ů�:�_��R��Ju�ֽÖE����K0��)������DLG.�ܻ�!"�#2����.������-Y��ƌ�a���aQ��8��G��l� t<2j*A�=�N��7�Jv[Y~����y �xSqn?��,Y�?f�\t�9�����:p��H8<�%��V&�j��B��'���$�I"�L�zB����2���-�ʔ�l|�44u�llB�J��7��>����0��^{vUB[������X\j�]#�ξ�/�I�`��s?�k�XwONa���ݦ�ee5x3Nq���/�.��od쎛EV��00
u�f�>�sY�2\�3p�<��7rF��k��XE? iP��A5���բ���F'���tX��VK|�ZD��s!��dB��We�w�^R�:���v��J:!T�P�HO〲�J9����	?6��d�����n�D�T�(F�H(׾��).ZF�::@���X�	U��R���`#1�XO�m�	>5wh�pg�1��~���։�{��I	#Gs�uf��.V�LTV�
s��+��!��t���|�# {�䢷�U��Ή|�qe�LxH{�1����|�$ ���w*�(��{��Q�����׮;����65��t]�1�fq����eq���~��1m��"�62��q���'^�d.�)�l�2l�G=�rXӇ��Jϡ�2�z6�Ex��tB�u�i�
��j��g�6�g��r]��y��s���3�[I��96otabhN��JѺ�s���ۓ���+�&4s}���&"P�w��iV�\U!��x�!-$��P�J��j/nwС�W���W$R���2�T���з����^D�{y��W��{���,x����,<}�%���8�I6�=�t�F���
��Y�,�q:U0Q��������� \P0�_�b���&E��ِO[#í�����>�xJ�_��-�᷑Pq�[�Mt�M{�����j<�L=,73]$C8�<�l�}�l��Q�_!����q�Ҧ�i]� ~�,�ʉ� ô���2�E�e%��6��ڌI���<�����{�.yd�,��a�w�f~5x��@�#-ʓ������~�K���=���a��NOF���4��8�`��64Rz���Q�gK��Xe�-��šQ;�֒�'�Dsj$x��+�u<)��f��#��pu\0���q�� ̌Ys�O���ϫg����?�	}i�S&[0�pPF��X�幁m�Ԓ�}�-��u]�8fТԯ��
`��O�45�DW��S	��ѵ�S�e�A�����Aa[ �3�(��P(!:1F�L�z�sｑ�P��,�� ��L��"S{�.Kb�Jyy�v�D�q��N�T�lF�#�����ҏ��?��8fkU���~�N0L��.8Au~5��~���y�h�A��5���W��Mӕ�%'������b�j5?�ղ�_�vT�=�
p�!�K ��p�?�AZ��i�maZ܏��� �.�ވ�i��S�σ#c�� ���X���9��p:��pr~!-�P��ז����T�+$��eiR�?�Ė����~�a`�w��`f%��i㠤X�f�xl��g��U��D�"��e��4%�h�,t��N��R#�W�	\��Q���,�z�;yG�DLr�:j-X k�`�)o��]8����a s�)� `��t�d�D��@�G��1ϥ��)��^&�!&$�'�X34���uU���5��lXV���`FV5bՉ�1~Ȩ�,m���/!����L}�	�۰��� hP ��H�6?�o�]�s䵦��u_#�cp�Ct��k��'?�l䢌ao�|fV����4���)dB��*5p��79�|C�sșsj��T�s�-mi{ҐQ�|DyN�5�g=K�SyI���B+�sJ��N��L���t\LЀ���Q�Y�ތ�� 6�@�Vݳ�DV�����/���X���!�?EN�͓���>W��S��6c�e��օ�?%�/� �ch-�/9況]��ʮ�)�l��$�) �R��ܤ�K�:}S�1Njb�W��,�*�(r8m����ɿIi�#Y�{!��w.XO(�!���2�E	H[��p��-[�{r3EP	=J�ͣ�31�U��|���2\1�_�ɶۍ� O׳͞�Q�(�CЕ��BW�t���f����m���$�ҵF`p$��vP4�+�ˉ�b��P��9}�T �P>߇Ọ>��$}�6��g/	%��'"�c�b��?1�&%Y!.'#���/��{��á`qؼI:of�Ն��h@h+A�sX�Z��ӣ�^�!$�#̫P27�W%�M`��^.�Vƿ�~5����Y�L����At�_Ϝ�\ag�樘 M�\�"$�B�i��W�oԲ��L*qx?���|���Yƥc�K��͖x�q�Ȇ�� V�1<���X�~��^u8��}v�7,�Q�� s$*������T�Y��,�b\-�
EC
�ϴ�:�U�+�&[p躵���.,�7��ٳ�o�uiaH�X���*op���-��G�X2<eD�fb��˝_a.�®TVn)L,��L ��3/:�����[i�%?)���3��J�:n��I��y�ۿ��6��c6Њ��DM��-��*H�lc�M{�!ce#}�MFn��z�+����k��m���:�x��C�e��F�3������~����OW[Z*m�����������o�BQ8R
��3������~�g<���!�bZu����̛:�h{̻Ķ��i /JY�bn����2w؏�����q%ќuҨ 6���S�QC�{,2F�:�F�����_����Hۑ���2Ö�V���`맹�ޮi�9���?��|�ⴄ������7FK(�_1u�͗�	(Z�3�cI�bo��$�T���ɯ�f������\�`A����'� ���fd��G��?��d�p<OW��}��pwMŸ�8d��+!��c^��Apjc�x�lY��I���V����NG��4��|����JG�V���D�U��	H=�u	C(���f�mrg�oE� ��x���!��܋�2U��zKV���Qq_*?t������V6[z�w�`9h�J�IC!�F7 E�G��4]�*b����C\���(ʜ��<�1z$��Io�����T(������ovx�G��pH�V3��[6��Lr|B�)�TY�۠'wapB<~O�p������>��y-o���(-xc!���gmOz��u��!b
p|c��[!��A`R�">�n�����O�;W�F2���|����.�E{ݓ^�X=���
OQ��ͭ���<v\c� B�[�։8�6D�k�&1博ХI� sq��!���:|��3U���4���
����7V�m����g��\��{GS�;,�{:�N���B�Ι��Yl�@�W�Wk������#����,�-Z>�x�9*��a�'�Q&�6
�L�@�On)$K�q�CJ312#ɻU�/`kYHQ@�`��,螺�"���N�z��y��T��P��ҭ}4�`P���s�O�,��#��w���{�L�#�(��֙Ǹ�w��'I.��E���6�E���\,PoρՓ�f�ﭤ�Г6��;��Q��&���~Bq����ߗ�`Y*�RN��R&�0��O���m�h�P,������w�졬��=��E^��}�wQ��{���W�3��	)���I�p��o��Sz�L�TO�|%]nO�t�|X��6�M���}���tH:��3$�:Ä�i����f�;�7�)�J;�Ђ��;2�<����l������[0��m;wղK^B��e�bKT�%�r���휡�aiz�> e?BA�ZU�e�;¶w�K�̷�;P�TZ�X=�{X�M�e_@�A�P� �?�5J9�eFv���b^�|`��ݿ��=/�� ����q�SJ�9E��	���5L��ReA�U$.���+��F�T�'+=|1-f� �8/d-�,�Z� �@BH6�5ǹ���� ��}~�����|j���C�R`�|�MGף�Kǭ�ɑG�G�_{��<{��Jf�޽}o1�ʑm�2&���d�hk1_~��v�"�"��;��u���-4M�o�uH���{���F��?�1�o�m�IE��V�\q�0}Ƭ²�wX��`�pk59��48�z��wܢ@�d40�j�l�%7��]g'j�
���g���[�Ex��j��x�~b	d����@����[�֗_�0e�`��X�k�F� ��O�0�Y1�/)����bd�A��6����Z��Ɵ�2{X��t9p������x9A}n_�a\�h�Z�;�C��D�6���^0�<c���]W�D�XBФ\��iQ��p� ymvg��i�m��/��?��c�i�ŹK�(<劀�g2務�±݄u�ɓbD?ǜЀYCr�َ����fW�>������'��Ն����r	iD�Ag�\�D	,��B�(~���M��
��we���W&�JKMm��.[�Ϩ����:�=sӍLIk&��!��0���E-%���q"�n���	|�:��3��7fڪ��U.�����g���Nr��(�Q�+Ψ?��	��� *��JMi�r��2@p!�r�/.�D�C����_H�;��S�$��3�&��TYg�9+��mI�AC�՜9(�����m�E�j潀hLQTG�B����ٮ���~��S{������	s:���:U"v��q���@��[�`�)��4�#�������}5���T	Q+�V+{},|�N^ �����8ԥ�����6X�H[s715G}zY�/�͗�Bk=��*A�f',<{���"��~��f���?����i�O����p��_Vjx��A�?��WFz�9JQJ��g�ZjKrK%���`�./F`��7�6��2����s��v�F����+}�
E����Jq���K�}#��֢Uʈ��ph�oN!(�%����:�#�<�2�*��o�I��\��kb�,ն"LY)Vɤ���;�|[t��9�t���t"!�0R/�c:�o Ƴ�H��34L �����21 �F.s�@%F�mK���TRL2HC�#�ቇ-�>P'G�zg��A�.f�+���*��2t%�D.�M��	�h�3R�DA��%�����V�s�u�
~�k*�xV�[�|@M�o��u=uϹ��e$��	y-�?���a2�uݸ��1"����7�c?��X��l�0���Z��*�U^�&��J<&�
9��D���t����)q�;zN���t�c�������R;5/xe��?
�rNѻ��p��;�����𵾑�e�\,t	�P4Q�{:�>Gt�G�7D�\r5���B"�Ԧ�n���c\�.!�s�Ʉ2�<��y؝�H|�*] 1(h�$�o����!șX�+��]9�����4UkS����PW9��E����`�$[��Ay�<%+�,X;��hf��ԏ�Q��%7�a�p���`�Z�ꞡ���o�S�0����ӻ����`��_����زSe)#��qȮُ�<������0�uΤ�Xg�_b3F��b~�di��k��D�Rx�)�r�^˼ˇ��3��M�(\*�տ?�Y�CT�ǒDL�m|ux7��,����yA5��0��hy�a������Y���զO/���������(��� jq[�bApI�M{Ž�4���Sǒm���U��k_-!�
�RP3-&RO�c�z�ޠ�D��)��Hqvݱ��+�k�>��o�B��۴ W�4�ב墔��Y��ޒ������*Ҋ����3:���:��0\�g�?�V��ۗ���ah"UY-Z(h�)�:�9y<-ۢ��;Ր������b�XV�x��{~���"�ƙ�C������yʹX$��	:-��#$ޮ��Il$�@� 
�@*��.��m3�6c|J_� Κ�9�,|9̐R,��?5�)���z�W��-�{�}ɡ_���G���e��^���K6����[s�u�A��W�{c�b��T�=-P�9\�t`����-a���9����}
��[�X:�(v�9Gb)�.޳@?M��<�����L�M�F��l'�^2��3��;b�ŜO×��,)�FҝW��?�Vz /���H
$���H��i?���׽���/(�
O2�7�xCs8�7 H�:}��j��7�c�~Y�+��p�m��Y�e���v+6�lP���z�5;��!�+Ec�:���	$̲�~�6P2�@�䎈 rU��"/�sASW�)}�uX&�	&!r�\��e v�2�^� �ڷ�ֲs��}Vz�@hϩ������i^
Vāy�����ea�v�W���l��{�8]�
�r��7|�U[!Qb��-REj��pnVO�x#�[f��Xy뗍��̚�o�4ahd��	b���)4e��+��PD�?:W��5�J���ph�R{?n!�CR�3C�V��^6x��ȷ�Q�g����u\]@Zb�t�L¸~b�?=Wyκ�(���{��������c�;���`��'�A5��C�ٲ�.�Tq�N̕}�Џ�hu��e_�o���,���»ܖ��l�|n���~ʿ௧K#I��u��V�݆"�E��Zjq�F���6^P�(��-#�t�d��p�H�K��uc9��<��3s���ƺA�I��管��1��6��#*��^�٥M������]n�-;q2��B��cx��\C�)�.{!>�����F9R���C8E��V�d�7h�����TC`"J�U�E����$����U��B�����lJ����5,�z���l�j�7v\�>�<�Is�qц�QJt':��+7z�5f_c{Qڴ��z6�����2z�EU+�k��qQ=��+獕����c�ǦSO��Xbinl]X/�Bt�Uu�W��J4�Od�ooq�	'f��^�.��גj5V�Y~�%]	���d.��t���3��(,��x�z����J��T��+%�+H��zJ�M���?�����&q$�yэŁ��ݖ�X|�^���En���
���>��.y�뇘���3�6���~3dA����;��0���f�V�`��71S�����3�S�(AT�����*,��'���~2��f��I�r�ch�jVV����uX^����m�!Y�d�دvp��W�,��]����5l��{���+.�!�0���Q]�_�AN#]��Lҟ%�zYn�u%�He\��myi����G@�D�~�+�};rupY�N���E5s�'��Q&m�e
�G�q[�w޽���ƃ}+f�[LT�C,���wN-�+��O�P�\R|�E��>����pkI���@�c��%	+�̝�^��]JV�s�uX
)�+Ԁ�B�m�p�Cmb��CrK1mUWh��SE����|��	��"LC5U�΍��D��o n��� �igL�N/7E☢6��+�-�H�վ��~��E�x,nfkT�������Ќ��wA�Vc�|���}�Gw?(J���)�~�~?��s�|�����q��Dg�:��O���V�S�#r^4���C>����\E����7��+⬑R��J��&�ۇO���p�P+,���E`fe_̒-���}�5�dcrv%��3�Z��`�Eu#�+�L��*�M��x��8�:	ӌ�K���,I�%�#�~�&��]���	�0�q��0P���O��-鏞A�	�*�8���/e����dV��+�/��B�~��<49&��3؜��ä:�N�$�a�������(�h�����+�	�zz2�С-
=W�~D�k�|��5N�6*2:��3�˵9����7@��a"���#�ة�IW�(�r)ygKV�g��jj����Ǭ҆�͎��=��E������6GW�̹�z���>��XPt5'�P�!g1cͩvp�6G����Sþ�����Tc1�#H�����m�� r$��PU���+��[d�_�4U��UGS!I)�( k�4�t�C��G�_�<�L���x�������1b)���!5H���ō�+��d��p]��xM�*��J�y(f��*� �=�q��"\r��Y*
�ޠ���]*v�ODm�[�U���6Cl$#0�;�ؓKG�W�sL`M[�1�$���3��N@��A�vy߇���%��]�	lGd�x��
L������FTU���	U�Éׄ�S��[h�u��`uW����	��������ǵ��l�Qa
��1긖��P�07*�������P���OK٫���z.H*�� �A��nM�m̧etC� �t,�#X'��)5�\� Q�e�t�E]�c��t:�l`(P�����.e��
J�N/�5nT��%���IS�@F�Br�@��J��,	J�>���?Ev	;-W	�j��[O*>m<1u>6�Î�K��*[K)A�&Nu�º�3j��g�@�����X�`��I�席�hs�>4�1`#�L�1���WT��`��d2���W�|I����jԭj�u��DT?2e�1LZG��v��,�NM�)�6r?q4ϱ�gP�JW;q�j8�2�������aP4�X0	"
,�d^80��o?��ZI�����̝�t'=jH����'fB�.ѭ�}��}�����WhD�Ϩ0���Ϊ�<%����	��,�� �-�*��)uۅ<4y~�|��F��Gq��Ia��t�U"&��n�����w���cڪBQ�2{Ij�~L5�qo��|_�BW���.,u��5߱R�L��^��$"F�����h�����u�L�Fl�l,��;��(x�!�;�Ly�o��E>�t��v)V"3�I�a@��D�+?���|sK 0��pwM�����ʷ�ٿW��ZҀ 	��E� �'���-.Hq��.Bt~FRH�e(�&ӭBi�ңC�;9�uᘉhT����BW�q_ٸ�9i�2�i&L�4��S�IA2�1��?�A�?S��+ɔQ��h&�ʀM����:���FFǨ�����Ь���|c���л�4/H�7��U<vq�9���T*1)g��Ԫ�>��=�Z�	z�w�D�����w��v��B%k�u�špٖ�W���B�@:��sN�.d \p��0j*z�I��OW{������n2lC���������@f@A�E��\z�9��zA<R!㌜�M=[����a�^�M���g���!:�O��-��Ý�׮�>�����8s��Fj�Ȭ�ss�K5��D�����Ń 8��Ջb`��&HSD��a(��	����7�͡G�#�	PoKg̈́�`Un
�1�S�QYLZO�r�55h}"��������#�G\2��XO��z8�W��7#���N析d9������4�hoa����%C�ψ��KL����r�f%��<�l~z.s#�u��]Z��~��z�.��,��/ރX�Xҷ4#��1R��fA���֗��c����șe�-t~��Ь�|^�o#L�m��R�^�1��5��𖨞�H���JD)٘٣�Դ<,���vV����p&�*����b��{��x%Ya�z��4b���~5�| c*�x��ɐ�{�~wW��?����� ��s�:K@�\D-5�*/;���~����LG���̳y�cx��&�D_�x/	�f�ܟ�B��Ixvh��y��%�?��6��k_�����Y�N�8`+�&�2Nl�V��0|An0َ�)�o��� M�1JF�-Ri�E������6TV��T

\�|��4���8!Ss����Z"C<�@<{��;��2�C����u,f}G[�s����d���+���?�ְe�,`��CW
k/oS+cY�H�PP�e��j��W��&\�\�}�:RD-�����;��1�]�<负(�\|�~h�B�y)�3o�{~�B�75��z��W����`�c�E��}��y`t��:�m�-SxS䩗��]-LfW�����Qj`EKj�������-CFu]-!v��j�38� 
��3m��>�"$���)��_�J� :��*G�|( ��%�^uz`�e��j������r�zqo����q�z���mbCҤ�,O��H��zW���J�u<��j��(��ϰ�>�i�d�b�Kx(�:�𲷎t����y9�~MU�[/rP���t{���5�0$�V��TMm+�[
��Z5u���xR�K��D&���W�.���:u9heB�уE[��?v�ϴ����4����,&����?qU�V�u��V,+��9'�FVf�$���'|=��_?�崉��!��,�]L��Q���,~� ����/})����r�-�u��lG� ��zx�]r.�p���fĹb�D,��ݟ��M�g�8D`X|����[�2J0NH���:��ZO����r�k���L
�� F�������dG��n�ՄLP��ҡ+֥�v������-�T܄>�>q�y�6��0�ՊG��0-����3Sz�t���9�g�;2���G�j���5Gh�6��ç�vp����<�)�r�ʖ-� ��3��t�����������bϒ�H2��۔�©�5�mf�`�
��F3U��@��P�N:h٨�z�7��b��Z�Q��쳛$�F�Τŝm�I�U�G�.�h�:(�%f'��ව�����束��7�����i5��z��K�!-��c"rV�B���N��շ�E���������j��\~�t
��)l_��v!������?r��l��-Șh���P�)?< �����l���˟��ja/P�,�G5+���=��3�E��<����H�;/�,�B`��Y��?�&��x�������~Z��^Ǥ��K�k �M��|�6���4�l��/�'�ӷ	�J�{��O��9�*��(ak&�W)3%!,kՉ�-WuѼg>��NH ��i/�g����<�R̨SO��ae"Aq�m�P�K��笪y�mib���ak�m���g~2�D}H�?����b��Br?S�j?��/J��C!N�-�7͞����b��3
�L��2���z��lG�ȳ�����F��\/_Q�]g��VD�L���!xv+���) @�=nVs���ߘ]�+�h�h���qG�,M �������v_ꥵsv�����YFV�9JF�Min\�����K�2{a�4�>4.	�X6�����b͇LNY��߯�q���fMؼ@���S�W�i�o� ���A]wM�,_/gi�d��KФ�S��:�0�:ˆ˭��-QX�|�g���D�X���Gr����%z�E��`A�c( �?�k�هq��n���������}}�t���ۏ�
�L;�Ձ'z%֭�J�%'��(���K����b�:V�
]��U!2��qB@���w�i�qSW,������p
��sƨ�mIn�z��ex#u1��h���0�"�&T�$�R��$�մ���1��3���c{�Z����T�5�S�D/��b5���7�b~Q5#��#=���f�4SQ������vRQN�Ū���6=b��.\�&1J�z�3�p�,Q��e?��j|�n�\�q�7�)�{�6$��b��c�{~�׷Qh�"���h��_�-c��#.��J�ш�T���n͡'�t,�i"���%��t�ؼr= ?�Ie^�S�C��$Aޣ�}l���+P{5z�^���	�"�2;�l9'+�\O��M64�?�]���J ��f� t�a�?�$����KE8�gn���"���;�Ʋ8��%����D�u����>�M}� $uq����npr]^v?^��� A�D�
��Fݯ��@D#�c?Y͋|Ӌ����!���<�Sf�9Eه��\bv���Hx�<O:�G��q�.mԹ����v4�ͼs<y�������?I-#�� Pr+����!�*6�58�A>��i��R4�΍����߾�v�ܽ�����ݫ��m��V[с�k�[�hW�@O0���ZeN��h���m�uiTq����*;�IWX�X#�Y�iw�wѡ(�E����W�YS%c Vk�E�7��涄��^M j2m�F&�IM�ߺF�h\�c���PCoyQK�j�c)��K�.��l=�Ș�p�q%��jV�����ا�f��<L�C"�f�O�9s�\��K����c�����=�ý.����"���|�s�9!bĻ,�%�/������/�\��P��]�{��K>P�m-I�o�ޭ�ai�I�EFZ)$�c��DMփ]�I!2F�B�;�p��� ug�8$��R�p�9�f����Ip���0��ʹ6"�P7�} �� �1F�{m�ብ��gU=�8V#t�ؙ4GվӒh}����3v���g��f������aJɚq�q�����v���T���M�7����r0Qg���±ڻ�Z��XUa���dDO�]�+��sLq-M���L����/��>[��(���������jUc��	qi|3��ԏn�}p}�9��{�b��w�@�A7������Z��m���Q���`vm2[�m�1Λ<1T~)( � r�nU�_�(��5���S�>�?�ga@�>��9����qFr�}�:	�b�Egn�SIݺCL
�����k'Bみ[#a?K�"�B�#%�(����8��M���CL:&iߐd�	� Y׉�6��)����f����(�`��F*�:�S�}���	`��!���*�Q޷N�����E���y���_�w��?����f$̆͑j�GϚ�����.���1�I�0�kS��'K�Ob&N��1�@�ȼ�	D�}��R!Y@����K��_g-sK_�����,�A�h5tY���KS>ۑ~���Ri}�_����xY�]hL������]�#nvz�ȫ
(�m9��Ĭ�����M�9�07L�S�>�������*��bsn� U_��>�ƵG3���H��˖O��W"��x"-ESX�7��`Ȗ^Q�f��ȆFc6�ֳ��.�hH���n�ϼU��;ڐ �yx@���2�_7/����M�u0Y�Еr�Ɲnȋ@4�%�9+��Q��
�{�� k|�j�0�I�M ��#Z����|޹�j'l^�U����%�L�%pI�'�tYёok1���/Rע^�X���������Àp�҉]R�'�iC2
XCQ��Ս��Y���[���yq�3�~�7��F��g�?pV�/k���Ք��ywb*'�+:��������3S���Q��6��UH�K�r�K$���O�n�˿�h�Q��b�t�"��!$�6Cy��:N�uC	k���X�Ȱ�?�&"5Z�H@�"4B;ؑ���#���06ἝfM:�[[D��ǾX��o�w�TV���H,�0�7yV&�}[82�?�7�9��S�hUA�m��\��V)/���j�ZO�m~e^�fߋ�:���Q��q�K�G�f��ٯ��9���Ơ�8�Ղ"�sl[Qǆb6g��+�w�j*ʢ���E������Swn<q�ԩJ�(�5�I�A`����2 ���k�-��A�Մ��>T�I�jǗ�\G�RBN�\)q�5�h��5�&t�`�`�-�vJ(ß&o.󇃡5�"�#-GD�vX��N�<�t[�j4eBJ�U���ٌ�s� �JDfT`����L��R-��(v���gg����wl�k����.�.�{�ma�-�!��o��4��+��p�+o��%׋�k�UzH�_vn��u'��礯���O����35�}qyf&37fa�2��\"�b���[� i��K�����oI�;r_����S�PL8{�E�t�ב@3�[�|��J/'�L��D����8#;�1���r��IM�'�/��B�����ZY�Rg׀�p��m1����}C�Kv�3l!j�W��K;,b��#Uݔ��jxtlM�p�O�yUX�ߍ���J9�t�}L,Q[��$]fF3p��L��!RC��;��u���1���,袚��� �Y=��rR0c ���Çχ1�8��-�&���[';��KZD�����1M'�!״�i�E� F��co
�aZ��L��Ң��rɱ
H������?�?@������#�}������� �:+~���+}6�(��l;d^rsfe:�?^/�9U�9��h��j^���pޏm��Y���D��;H�j^��Y��T7'�zhY���sa�`��<ύ80?����=���V����5�`�#'H���`����\J"R?R�s@*�-1������>,ʮX�m:�}_0J7�с�i��?��drq�$��}'�u'!m�����|��8�o	=��vr9t�>eNWlƂ|��f��\�U�ox�n�:1���(&0V�E��I����Y_`8"J��s{6��P�CW_R'=	��>ޑ^n��!�����Ӧ"$S��U��:0��Smz�V�#ywY� �N�(���<��[6�5�����ņ:paB�AZp�j��]e��%O��"鐐�2tCT�L����s��@⊐�!���3\�a/V,˔~��T���H���r-}FiڷK��j����%5�
D<�Z��U|�P�BX2C#j���i���K�( ��#�T�>�-�JۡȔQ#�f��T+C�����|^!����ҏP�s�쒟r�S��;�4+W�o������[��~��S����o�̼,f�B��#i,?? ����x	M�f�4Y2� ��A即�aP�'̔�>�[�]��C1M`�T³b�ۖ*��_i�N���~d��ZxLD/}Q!Q�xhOloY^7?����X!��;�$�@�5�~�F�b�B����_c�>�c/�f�KlY�\�-��l�z����΅5bN��TI�S��'84�����?b�7��fyHF�k
��tb	�.F.N=CX��Rl��Fc�kƨ�����0�P��	C��)�A�t�j�yW$�R�Iqq�i���;s!x����w�¬*͓�J[@ƙ輴 -��mvQnS
æ�_Źij�13�<�ㆻQ�j+������X�(!�5D�/��o�)���o.���弬J-����s�`T襣��h
�:���^ �)�
i��VJ�yp�
�C�F?����VS�Ĕ�]�Y�����8J��Tk�)U |N��\�Z#&Y�X�8�tQ��`�Y2�tT����SmУO�(�`�_�\��%�`Vu48?�E#�P��5��, h<X�R�)�<��l�&���a.PeP=,�%U#�W�e�伇����=�⋧*TH�{�t���t4$P���
���+�ы�[��~KBc�"<�Z�'�����s�br�Vk&�X^!q�`\��mE�ǜ R1!�Gf�X_�&��zo)���4�%e
��	�m�C�B�i�t��EY�h�ou�n��9wX��4��xE0;��2����+H���L9!-� y���7B���C�wvXW�\ S�*,6t��g8tC9$,^Y�Tp�X��e(���Δ>�����4��\n�oԀ ���r��m�uM9C��aa\�I9E<��H��������JW���~����g���-9
׸OyUpW�7��)���nD�w���F��C�m��f�S��cd�:S�5�Zlb.�R�3�����wM�򴷃���� b�F"Bm��巛�_�����oA�l�[���p�B�" #���tOܹX��)��qh�h	4�ԀVPm�l���;)��W
�r;=��X���QA@��:L�J��VI`�Z0���B�s�#�[���2��S0�G ��� ܸ��C?uC������G<��)>Ԉ���#�yΗ  P�Rf�$��[�H�CU��j1�˨`���@�8��m>�+\I�f�v5mI����b1x5�嬋�D��Z���Og5ύ�����g?�g�E���P~sa:��&�7z6�W�*���ڻ۵���$I�?.6�:�X�M�w��-�ZV9gԖX���ŭ�s	��Ǣ�Fd2Q3��Ga�����~�5�X�5�)��2���0����m��E���.(h�tG�A^u��^��D@�(.��R��D�Fܚ?b��X7��)4_�}� ��������y}rjɶ��#�Z?��`0���@%�V�4���ܞ��5����Q�p�n���~8X�[��Y����f��MS���z�L��.��:���S�/�rm}�����-%�zI�HQ~S��E�d[:�zKO�����{a�s80e��K��+�b�N��l���{������Y�W��i"⬁.c9&���ۼ@\~[1'Qm۔<��Ȟ�t�\:CZk��{��Rn���C��YE&_���$}�Qݨ]ӫび.��Zޤ��nkƙ�I�Q<2�W�8&�ѽ/��ݔ����z.�26��0���P�ez�J�Ĺy���uW��5r�A���S�-A��@U�hQ����آcpQT�V�`�:� lf��)+xǰ�R�Q�H]6��2�;_�-�)�(�ۈW�IO��
��>��?a{��d�o�Sq�ڬ�B���*5r�o�Y"��_+F��4/V>E�5�r�4i�5&רE�\�qK��k������<�SO�N ����l�Ҋ@��$��Pl!!��9�y!M�����f�lY"���pP����6n��ք���-����ٌT'�'�P$|W��Q���\W��cS����Z1�a`��:�/0̯A9����v�����ʅQ9��!��[L�Xd��3����C� �;��������������^���0q�7�����*�ԑ��I$b~>,+��9��HCO<�~�9��q�&�Y�� +d���^X@=�R-��{�rW��mo�5O���IXQ�p�Z��c9}�vH{����"Z�
��w���,-�X	��m�*�5 ��~T.�꥙X�c��������V	���& �XFk*��$a�z��Ű�W��4��g��E�0I4.9Q�N�>]�a��4�^���v眡Q(&V�9�¡gÌ8���:���������~���T�&�n�o�а��g���f����?S�+WF�;V��>+���*��5�d�|�
�t��=m扤�� �k�y�_��+P$�7uB��Vc�jh��/���|k���e}m.��j�`�I�4k�򈰬2^��]eާ�ģ��@Ob��r��)<�Ck����]R�mC���c#��t��|+7��I��~O|��:��P������� _w���<��n%m@GL@n����~uU���#)��9�>N��R���(��T���7K�#=��Lk���91����?3O�*<fR��fe-|�;ՈA����	#�]I �g�{㮔����a`�����$+�	.�qp0,��5��I�w{I�0N�>tȥ�^������8�\S���i���|c/������=���p�j y[O�л�����ܗ����Q�M�����ضc�~G�d�jS@�y�-
-�q� Q�B�P>��������e%��2�������Y�m�_E���}x�ۂ�?i��}�Y�#�=�����ߑф��Ŷ�;�(�S	���E��|�8ߛ��j�Y����;Wkb+pM��Kv��+�B�\�����э�ѷ��Zb�7���i	Tb>�G����'�/�7�<1�z�W�z��j)a_Ԏ�xi�2d����Vq�=�D��q2�t���V��^%�X�Vѹ>O�8��G_�͉o�p�Z%_��u��s��C �Pf7?i?���&	���T���3WY�C��w��͝#�"�|F���Ŀ�gZ:#�p 3%��^5U���k?p�JlfB�Sy��ܾ(G#
]�a���5Pn��˨}������L�3���p
o� Ϥ�
7GOR�s3�3^�V@I��)T����9���܋�L��3�ǃo�-��G�4�c�U���D�,�L�}g/�{X撮�����p�.��$�"�W��g��1ώL_��XG����YIb��Z9�}Q����53%���R�a�	�ƞ��M܅�hw��ujȋ�A���Lc'�dv���2|�TҸ&_�$��T�d�A �n���8��$�F-7#Sta$T9��R�L �/�Z�H#ŗ��?�.3o�Y��˰��'���M.{��{�v������"J�&��׶��R��/0�D�̛HrtLYP�GV��� �r���J5b�0�0ȃ��]����N_�2���U�����N	q�g{cN����;`K?��W��N=ϛOp�h�;�:����/a_�B��(|������8�������e诰KY�O���/<C�y��˪A��UNy�����<|��JP&���Z1e��ϔ�rs��ѽ|��?��Y^��[�2(B�+e�/�m&$�d��]���7��C0��� YR�~���T����R7U�<�p3��zb�,�>"�v������$8lb���>ڔ)�f�}�1�éV3U�`��U�h�^D�zA�-�E\�H^��5�b�bK�����âW�J�N�~��)N9%E���EԤ%mT�v�e�M$��;<�"���kW���h"�uɴ?W���Zmν���^Η:_�C	��?@��t˒̓{ʋR����.X�Û(:gǖ��9y�i��9�
�sN��z��JI����˵�-&�g�J�[_�N�0}M�[Ջ�ת��2���(߃oڱ{j-�3&��E���R����pJ5TX���0- �'�kSGܺ��J:�]I>FM���S;�����v�b����5�fl�������Lw���^��b��۶�Z�+���{�R���ǣ	"$���Yx�F��ꄅ^[��iD��3#<LfN�^�|=�}2�:h�*�
ގ�Q��]�/E�.!��6(I�m�}9��\9"�_�32/�Z�8|�12�b�|��5��!��.9b��M\j�D랻��j���@~��I���c�l�[�����5�IS�μ���9������8y��T�r"�]?@Z��H�s�,���iMm�mT��F+@p�1�Л�U�[o$�9=��������Pľ���n]�8������Va���A�7y�2�Z�v�J�&0���'j1�m��(��8��{/��b�Eu��*�*��&=Qў鯸��Alo��x�<�)��h��<7�I�.��k5�]r.�T�bT���d��z��L��� ��[xc5��R�x�o��(�F�=x -e��5�s��~0���[s8��A���V;=��Y2������xkI60�<otG��z��H��B�V�r#\N����+F���H�lv�=|n��#���Iѕ�d���c�����T6�΢�[FuУ�<T����>��M��Gt<�͝Jz�d���k�&O*ط�+v��ۨ~��)����R���D�_�� =1�91�n�V�y�B?�kPS�gG�����3���ER(,���HS��r�se�=�k���v�?� ��K��;o8�ּ��{N��Vw7&�-��q��~�w����'ޏ�mY�6h�nX³���=ZEc�j�/U�Uҕ_���D�_���u+��8I��`�Mp������*��x�2�3�����P{��	��X���r�|��D$����͌i���)��LS5����v��F�-i�~�j� v}��=�ZP�#雺Ζ���
�TY�e�,���t�`ڛ����Q�� �.%v#7��$X�N�A�r�T�"�u�$���f�h�V\�C��>s� a߉�v���yV���m�g�fɠN�ۆ�ɬ��~�<��K-U�~���R�@�.��h��a�as;0m�)���6v��枏@{��>a<����p|�	>���XOs��\�&��O�w�i��U+�I�N�/�
��DQN�{�.��8��Ck瞺��&�ᠴ��o'ȝ)���Ey)zs�p��ٸ$lsy�.��������kd�$2�$���o�H�A%����0��,���h�%[1�d�30�^?Y {�P�a��ȡ����sl �U�u^.!�p1I�E���}�=�5��[yg��B�Z�ݎ{�������n��5��y~��36""�9g�1�v9��?b|�k�I�[�@�"��Uȡ�N�R4e�b��)��+jk�G��jѴ�����gw���x$��$��m�2W�<�k�,c���C��������E�Ƃ�=/;L|)s�k1[Z�@Z���L:�N��]�etM�YD��Ac��^x%-�ن�Y�F�n]f3qh���O��*�c����;V��{XiL��	��Ri	g�0�M���/8�ސK�lKV\)�>CP��ʤw�0����r�5)ȁ��(�KΖg(�P�����.���wخS��͖n���U���;l�B�����J�b��B� ��[-�1���Mc6���} �o�@X�ZJ<�Imj�X�[K�����ONQ�p���gɬ�C��!�;5*xZ¯�³�x�i�,�J�^?����9�,{]s�cֿ�J�B��o��`:�ul�b�;2ogOS�1�3�:�X}?"N-9�S�5���M�`bW�����gġ*3���g��/9g%r��
I��9�c��8_��W��Z��Q%"���d(��aѼ��N���8���"�I5���+����Y�z��{hJ9`���S� ��F��eo��*��b_���Ĥ�_ni�afgfy��.G�P��F#�ՎC#�EN�\'�B��(�Z��:C&�
�"���w��i����o�=����f΄r�in�7�ȷf����0;�`�s��,�?�>a�!�����-�M&�ԓ*<�!h$���N����G}(9:�݆0�	�!�&����m�JҤz+������q!���L�N�֔���yx�&�~��o��U�6Rl/[կd�c�ë��=غ($��e#��Da)o��r��Z��} ��K�]
��:}��AWtM\�<K�r1I+ QR8�6�����>�:���GG���޿S�O���[E��d��xB���7�����0�6�S��m�{�i�~�hj���s��Ĥ���`:��LC�[$,!�η�F��9o�䰕e�J�w! ��\V�e���Uk�<�$��5ܨ%u�=�&Q^�6(�O�S��=����t����ީ�]Lq(�)%��W���'��"�K�����	6l�Ľٮ�q�;��(��\�~#�ј_��|=%£*��o��64�\���=~�l��������m:t�Z�n+X�0�k�B���}ܱ���4`m�*K+|
���q0�K����IT�t�~�i����6B�f��j;G1S��]��M(0G����{Z�oHU$��=6����b���{�����'B�̩{c6��g�`	���M��0���Xw��e��y��oX<��Z��+��?Ĭ�ȶ�K��.I���_�Ϛ�縰�Gz{�=��IH�S���Xn�ի��ɰ�k��Ȩ�fN	0��(I� �#?|ß��H�p�4����l~2�af�C��,N�L6m�s�#*��i�;r�[y�w�%�}x���A8Zd �{^˘��N`	,Υ���2hO~�mKr��T��lg��N�#/I�XWё^N�sw�ɬy����O��	WNK� ha�V:�n���L�;� �0���3�7���c}�ݟ�A�'�an�;Qe�a��N���u����&��-* v��'�1Ih��u��o性�,*}���y��T�>�8�Pӄ/S��`���1/��s���4�	 �e"ٮ!�M��7�i)0�;�E1OR6���Ŵ��7c���A�,���%1�:$��]B�	&�2�P �A~b�S:�QDM~g������@\����������w4�vN��n\���Y]`�� ?��!I�w�̥-(��Yↂ����+Q>K�>���K��h'_<��%nD)�����/rS����{�*x�����̤���[����������7��e[�;~ٮ���aM�f|3���ۂ>�V��zsvY�6�����y�rV>g�̓2��״�vcנ����b�F��bgz�F*��ō>���0ӕi]X~�Q���C5�_Ǒ�?�\!ڄ���o�4Z�Wb���R��T���O\ b�z��
��]�Ĺu�4^-�ٴ�]{P�k8�S�y����f�GBnW���/d�09�0�V4|\�|B����Oo���"�F����_v����J@����(��2]T��n�R�48Oi�|�£ZHT����D	`]���>�n02���t��^i�f�+�Q�Ж6ݢ_	!۪3��=�wHJ�[�?+�xSHu;��3�;JR"�6�0y䱪�{6DP�qyaI缔^����H�>�;�v�٭�W�-�S�L�k��Ӭ'���nk��V\E�h~;B�����h#���,~��xF�屫-�z�J�U��V� �?K�|��W�;J����%�S���?��R(V��Ї���D:�Asوs�/�{������ �8��D�1j�7ap(/%�-�����pr<ߗgD�n��G�g�>|T����Κ��	��t���bL��!~�d�~������5����G3f�,dWw��>��n���=���5�����ݐAS�:�μH�-O�7��ǌl&��Ц�^_�D}|���؜�V�i��o�y�3²R��_�i
����E�rA_ָ�������ʥi�*څ�X�웜�&[�=�3������6��z�mYV����a�;*B�������	l�B���YR�#k��8�#om���S�,v�k;Fs�jd��v�Ѵ�H�#��Vp�
n21Rp7{����}£_���l򴳅�KGmO	�vr��r�ģ�E8���t�1p�A�'�/ر����h��$G�!^}6�^��e�����������������w�L�5ԀnzEm�C���1	t�Ձ��]��' � ���	�??��ɼ;�^�Ζ��3T�*���$0� �0ꄨ~O)+D� �!lԪY����k���.pu��"f�({�l�N 7	� �-&�0�r7Y�׼++�9��s%�ܴg �E|L%��Sk���3�7����Zls��sX��	�u�I3F�'gy0R�Β�?�w�����6�{����G�[����T�_�ȣ�ȕf�^#eN��O(>�MF�o
UY�
��>�5��ϩf�����B�Ѵ.C&{Iӝ�G�\۰I�
z?}k�����!i�;���G/.�DHJЍ��$���[j;�E5�=3`mŖ��/s�+��I�`�bwѻ�ᄠ�i���^�i�,̪O����B'6��G����ڹg1�<)a������U�r��i^�O7�	�ev���TV��ڗR5Z�X�9�<i������<��x���Kk{�_���8u���P>K�fP�#�IDWk�_��L���c�ٕY���;݂�AE��G;M�Rf1�=��}�j/n��z0Z�=f�(����v`R��c�� ��T��y��+��|��8���Ӟ_�7t���4��i�����D�f�����H�0�+����|E{X_\�o�9C�5�A��UVRNQ�D�F3An寯ȮS�lz°u�4~C���8���
�@
`����Gm��W�uB6ktw?LA;�t1���v@��D:^/ؽ�yor��yf�?@���ג�����P�G�ܡ��ǀ��JX�޴��
��}�IݣV�k�&��@�;�W`�B��TAb�dy]��X2��=*B��@1vU1��i����j�O���9�	-:��|cΑr�(N������(��Zq�,il�K��4+n6�R��!�6u}jO������QCa����������'PW0�[�?�t��}S2�8_R�E�ɺ7�W�p�N}^��%ˏdit��П�m��R��J����?X�?�z^��d!
��U���pbsE��+��t~S� 	��p-r	��4
����Mnܒ�;���%;V����؟�� ŅC�d�<I��y�;����RR�z�M�
%�b}6�0�ݝ9>��Ț�k�	gBM����R<N'�`_��p53���9A͇$����U�|�0sE�(p��L!�=�|�/����D�ܺOW��XJry�������d��L�b�B�ρ)����'���O����9q)|r xo�l�XvA�|��#!d���#Ϣ!8,��뵱�Y;��#U���s�A,�	�cx4��*������Y/[AP��I�;8�������z_�_�m|��C�6�y�a(�<��CI�3W97�9iAiHC�Kg������r���a��<�hc�=�D�|vo&�?/����&%�$`�dl�H�#������0$kkͿ�¨����z������Bj������i�.��c�їk}��}&s{E?�rP�&�~x]v|Yf^��u��b��.y���q:�Ba��Z�4���q�O��.B���9,4�إ:������=��׳��1[,�޳t��e����%"��:�p19A�PD������A��u�@��p�|��P�,�����Ncg�QA�ivE�+�@,��L/�0���h�"��4ex�@6��|9�C�4u��#ߝ���_��M�qS}&n]F���&� �3��-c���R����5�;��a$��C�C�q:A��X��"[S�i<t��d�d�9���.�.��?U����`�_B=+�����+�(G�#S�h����`���ؘ����,���ź�x����z�F��MH�Pg��b������T7s����Үr���GԎ̃�:���9��"j@;Jl=�����!F
�NxY8*!5z�zֲ�S�+ڐ����ʅ7W#lT˦�k	��*3]"�נ��̛/��M�� "~���lr�I��uYd�2FP�/��T\�|�1h)]DP�P�����g�F�n��࡟ZDk�P���M�}����J���R:k=��s��\)d�;pڡ�,y�yP]�z�TF�m� �I����]���/�||���sb-Xj�<�<n1�f��~Y>��*��ѵ"l�_#~�"mP=���{~�X�L��]�
�V�^�%�����!B2\5�8�����`�羑u�O!�aWm*���rUem�Z"��1����T�]�C�ɚX��+�ۘ[�1I������ܷiN>]���>��	qj �Q�R�l"j��(1��������ƒ
�k��������)`� h�\UفQ����f"ӊ������y��<.`���E�N�鶦!���.HiY���Yz ��D������y����7�P\�Z\L��y��#`���<vQg�4ߙ�S~G�=G��*����Az+���2Kն+�΁be��!�~�e^O���r@�{Qs��a���>:Ť�2@�j��b�\@hߚaޡE�|�:s��H�˲�j�l i[�jg{�!G�da�,��J�����;1&����/#>���[��[{���dp�!�q)�5Z{��e ݫ�0C�!Vw��F�{��3K	�����L~el�l��-�B[��S��!۱x;�%#)eL'��o�qx9�lf*&��7�����a)ZZTCq%.�'�%еXm �8��N�Բ�������M�A�aW�1}<�!��SCQq�A��Kz�i�#p(Nb�,H�M\_��8��͝$ �IgIO���p��v�S�+k}VȤ?��!y���R4#eT���<��?�Y��Y��>.�\�*��k��B�U�L
Ug�""gZ#�+�]����߳�4��>�v���D}���g��k�Y);�Q�6B��{*�2���?M�%���h�Y�H{��!x�tP�.�[d�<�ӞA	�L�:/'��,����r��<'�<�B���i�~~�+�V����E�,���E��F����C8o�(D�E&,��\�M�<��%�e��O9���N,L����٧�)DǄMT��/l��������^���'�W�<i]����>�u�Z�7��2`�V�x���Z۳~�o�O��Qϣ�1��\�D�qd��Z�}��_���>��a�JiKg���8R)����/��J�:&�Rk� v��v����U�nS�LG�4�Rb���ySB�}&����&�C%�c��^i^�ԟ�����Q� +G,~���M�Y���ʙ^�y���6��2�,)S����ZnX�Z��*�K�ΐt,�r�.��Y�4;$�ea�����:�C6�
��S+��*��y��>���K�7#�r�W��u<c���� 3���x�^�cD��T���l�K��"5�*t^�/�ͽ]$j�
�${*���8s�.۬�����:t*A���Idl���ȖU[�m@�*���� ��" ū�AltQ@a�2�bv�/���x߽o����M�b���g�0T�_���$��v�D�)��G�%�ya�N_v���Tr~�ɑ��;5��o`i���#���;�6i]���FW�%�p��ś ��y�zZ����tv�����s^.� ׌]Jo�vv=���4��b*���/T�b3F����H^+
�*���0	W�N�,=��ݐj�p-!��v�x�J�~&���h/0����d4���Xŕ.�ѧ�>�-�������J����)n��×�n�'bE�v��U|aM���z�,ͫC��(m%P�"�l�l��*Rh&ut2�?GvN�;�����J�+�_J�fɧL����Ջ�<5,گE�����h��+m�/�i�5ٳ;�􂂒]乕�J���aӕ*+��e�3J��>�qn��vY^sW�\;�\]����㰫}|�϶��X�@��[��x���U�C�睠P��W2��?9v�4�SW���ԙp=2 y���Js2���B^�+�v+��'&�C"�<6�$��d��	��`���\��PNi7+�y�J��c�Ȓ�k��2�
�!�5F�*�\��p�m���,cQw�����k��.`����1�q{W^�"Nߍ.E�"���E0��"�=���C�(Ct�kG�F��8���'/�+^�W�`?����-��1h��} ���O\1�Ѱ6��,>������olt�ω�%�}����W������.%��d[[���θA2)����f�dĿ+zN1_`#�E�BZ��تԮsq"K3Li�vZ�{���it��`T�d�T�N���lB�ўDdf/q"��N���׎(o1�d��'8�r���<C�3��*�E���>@�W|l����F�}L��l�k�`&�^��p���;	�/Z���� _۩�4 ��F�v����A�C�wn����Ol��f����z(�FQQ� ;�P�U:�`|��r�u�c3�.�z�9�Q=��%չ+�K��)Ԋ�PV_��y2�{J&���|X�b�~E��� Qŧg���w�3��hTK��S�r�ܡHq�����qڨ��
�5���{ӵE��DP��:O#D���呦������W�3M`�%٢���V���Ӏ�5<�Ai~�X1��nG]�/Z���3&�Q�B����m��f�s|���cş�aaMU��p�K�d�w�P���F,���:��{��"ou�N���MV��{ܞښ�H>��m�?򄸕lKӄ�P��<��q��$\:�n#Y;�������2� ��Z���S$�q#h�ϸ�۹4v�w����U@`���l.�.u)�Y�Q:�=^&�k�P�h��M��}�#I�ot�{�݁֗�Y~�x���"����?���
�@)n�цW�0S�c����������ɟծw�á�;�T�Z_SȜ@p#�Y9p69��4���7�s�F5��u$�_^����NKY=�율&r�
<�;�].(%e����w�R-7��0%��xv��Rvw,�M�#ٚ�(�Q�-�z�Zx�S_��wa&�9���<��YD�HWAKd#�iZ��B��������3���v���e�0f�	D���2��lu}�J
L�I8[�%dRۆ���a��RqP��SC�#��c�9QL
����{J�"�S�^���0�9������*�������q�|	h](H�"�ΞǮ�K����#l�YX�v�9�'�"\�OB��B�o&�|�8�a��~B�Ɇ�Y������5����8m7 X�v衍i*Z`�L{�Jcº~���[�P�AGa#�P|�W�/d��T��FU��	^o���|g1��?-t��60!i!�q��IB����Lm��)�+�z������`f�R%��T��CH8�d$��Sa�lc<���1 ߐ�>ʉf�[���,*�OF�>O%$=�-A+������w"�A� �a�jXtT{�qU :[��eS}�_�G=�L����a�h4u�\�G�nB-��hᵒD�ƕW��d9��+}4ɧ'�j���(J��쁌��W;��oF� �������8Ty_�ٻY=�z��m#��OZ�~�!ɾt}�u�]nC���SGm��D"6�T0:���y��Ɨ�+���mWk�G�k���5���0�p �c�Hr1	ba�=���a&���ʊ��@#��K�(�ky5�y}Bj{��m��4�ߘ=V��閾)xv���g��qz���7�)��tA)_M;�ҙpX:��j�<���ޜ�ŏ@f�|KH�s��u ��ޖ��~}F���7�{y��p6�JW��yr�����Q�=��i��O %�ȉmda��ʞV>O<�>���L&��h�~ۻ߄j�R��$ql��4�L������̩���w�WC�!�����OhFM�T)�S�;s�o�,�Gn��åT
m�$�j  T��� �@'�d���(xpi$��M�T6��÷қ=�>������!��T���_���߻���T(���%�Yd���Bx�^�0������N����
���i`v�OsE�G�>�[yM��F�7%�r�x�6.��������g�� Uy���n����,YIl�36���(Dvi�b�|��OM\:g�[j�4���,�Q����j`/�>=�n0���>�|�=b;�Ǻ�q3m�ϑwr�6FzH�O�y�y#b���~��*���v�Wc��V)j21	��B|$h�l�;�hZHmB�o����[�c�>Je H���?ϲa�?_�g����D�h��T8��{	�
����Mu��7�䞈i����� vG�r�0+(���HwI�7,m���ׁa� u:�;ǐ�JOC���~�����`t���т��O!����խ;]*��K�Skύ�|�B	v�>�j�6A��"���pD$7��r�����{��6��m%!l��H{����-<����8�:X;��J�w0V50#�4��%� �sh�aqA��l)d��x,�bK_A` Z��C�?�?�\�{�L�܇R�i�+wܲ��>���Z�c��"��F�j�V�z.�ok�g`b�7����Ŵˢ���'���(42�poMɂHT��y/O�MO��Ȇ���k�x�!���p�đ!�a��z"0n~A�o�v�(�@S���D�V���I�;��}e�T�޷�Dǒlr<b��T�z��C�8p#㒦eЇ�����Kl3���#h[�pu�w�`v��tr�l��BMC%{L�X�۩�`έ�v�+���Es�|��]�Ƈ���M�G�6	}{Z�,���sV>�oul�<a��{7}	�K�L$���h���Q{����G���L�\�u_&�t�+<#�7nX�+4r��e���v��Bi{e Ê�/��(gI����	�@�FV���5њo�2	'8�Uz��{���/�m�ݟ�]92`�)`��9Q��;L��~-Ʊ�-��b1�Db*i�
��S�r�@�/$��,��༭x�/%	:���̀^�D�Lc�������5.	P��_U��|OO	�7���#�[��g���<�UĤY�mQ�a��ȫV='X�a�"��q�Bv����i�v��EQ���ۉ��7X��O�;�J �m�X�nX���=�c���3lm��j)��1n�w4�7���{p O/��G����R��.T-�I��Q@�G�y��?�qDڻm�ə#!���ܱx�^?����f�E���MM`�$�Ҍ0����g<�4��ݾ[L���m癶U�[��z~�/�1:q�tT3v���u_���X��$ 6Zl�C{��)u��N3I\^F�%��GG8G���� j����D�v���Yn���}r�.��Jit��a����ruh���O�M�"���[H�O �e�-���0��P:�l�~�pT�x��y�N��Y�A
�@/�<Lrvj.Y�Q�xI�  3������SZz�r�ȫ�9����֠N�q�=��k50h�r�=�J]Z�PQ��7J�|�Ʀ� /�� ϕ��5}q}f��@�须UW�V?�\ᒱ%ժ�
���\�H�Σ>9�i����D@�j���!$O�rA�ղ�z�� �9��C�e�*��M�	�͆�'�*rwL��	z~�H����;��~0�W���ok��(��FAB��1���6���p}��75C�ئ��I��&- �����}w��F��rP&WL���Px�n���ד���;��e�������P0��/���=t��˪K��㯌=����;W�@H���औ@���4�w�Ͳ:$鋍����P�I�kkaV� �_�P��f$T�'u���Vit��f��k,����[m�aiSfK�0��Zs���1!��Sg7����1�E|�����8^�
O�[C���|��K�D:poa�YA��S�����*�S����j�Nڝc3��T�P~�~�Å��X��w�|-t�6 YT<���nv�n��hL��I}h�dv�6���5(��R��(�O��g���e7����?�����պ1iQ[<���!�m�Z�`���j�{f��b�7�3�;	F�ߙ[B�eI,ֳ���e����9	��0��DF�f�^$��r����.��U�!����j^��:�7��Q��䌒[p�v� ��
ƫ�J�$�U�G +�1Gh����I�K^�"I�H�-��?���&���	�b�I�_����|9#��:�d&��8��%2�jX5)0���C	����*L�:�_!�딤P8�.X_�7R]gH5�n� ��Wx,�2ݴy��Lu������|6��.$�ܡ�b2l`��q(%��WX��F��-e��~@�|�����Ǚ8�� �7��A����Ś�տ��԰�z�%�+�ec�i�Z��R�q �,7Sֹ� ��T�Tέ�t!�����e�߄�p}���i��5��J@����"���J�K�sY�5J"��r)�iK�(}���a��o��\�N[L��l��i׷+���RWz�}@Tt�d>��ͷ/
a��_�cC.�T�JĪ�?&u�%�c�V8��ka���>B�-9�����M M�͋�ax�0;��Xw�"�=)���į��D�<H���� ��+�록�=:*�o����������Pn��0�{L%p1�!�U��͋�ذp��`p�YRy�3AJ����B�"9xli��'[(���K/D�m{o�eQx/#��Ϧ��v8�w91��Z�A����J�t$��
sHe8(�օc��gvlC���^���(]�U�^�a����i�&�6º�?��ks���t��|�ܠ9w�9>i@�qo��qWj �i�+62���1R
��!��[����N2<�����H� āS� �)��b�P7t�B�`#��q��蓻m�dQ ��t�ܷ����I�>�m`��K-lטD���]c�,'9(��j�~B�R��� 0�:�n�S.��#�+��*���U�:�~]��>Ľ�$e A86m���"��������}U��M�id�y��伵�a�v�0�O�W��F������A>Xܳ�a�-X�"��*B-��@#%��80�{l��x�Knu�m���<���˙&ѲH,������v`��T-r|��H���=#�0�>��Zk�Xw�io�B`�2[�1U��9Sҗ�� J���/�Ҋ�!��_�錡�<��}������~Ԛ H�5I�T�s�L��Q̕(�V��iT�6�'HF����.N��_�s���#��A5��@��]DY�}'�뽓H�X�QM	g�R$ �K^W[�c�d���r���v 쿉�%����+g�M�`�������u��$���@å�6Xt���s�.Y�[�>[H����������7c�<^��c:���)��V��y}�0�Q��fM}����-(�n}���6!%��|��-ݘ�D�8^2o��e,Mf�Qӏi��rCb8���{j�ԛ1��w�4�� d�����%y���ńrJ��ē?���N"u�a��L��?���*&�Qy\���QX��k7N2������uxu��I��N#�AFE�iP�J+/���� ZPx��F�W�����$k��[>}`�1t��$�9����4%;����s����<׼U �k$���������T��.���4o�n/y|z�e���"�Z�Ub4�(�����<~���ܮ3]R�^E:�|�|�b�r_�;����@�q{��I��U�W���h� �����rv���B�
��駰��_d�221�Оi���񆔾�υXƧ�Uz�J/����+M�����ЂZ��r�5ұɪ� �-�[Z�-�#Q�40�)�����T��eYM�.@H�����������tID��L����.ҵ;�_O���ko�lN��e�lA"Ƿ���5B�˥S���0P�A�d�$�����M�C� Eh���6B+�N޲����P�i��/ ���
=C�|A��C�\�^�rI�ٷ�α��՛٥=U"ߡ�g�+]s)�m���Ht�-#������Sf@��/� p_C>/�Y�����b�D/K���羷���q�~.���s�Z|�&:��0�LZ+�=>U��[Vl�4�9�i!��$9�$��]w�V��!Ϥ-��D5BK�r�ɸnoЏ�+kg+���O����ŝ���߃���o<1 B�����"�x�`~���v�,Gs�ݻ�܈������������3}���R����gzfn����N�_��
�n��暓��-W:�wa�n����{Ȟ�kV_��z�v�&�U@��roY!׫cNw���9������^1Vw�����	cp��|{5�w�ZH�u(�^#�&���<T�%�g�μp�˭[�.�6�XT~=;1%f�y#�;j�R0)�����I[׫�*rh�G5v-�����)"�h�˧�$D�m!�ú+�����g�o���w�npC��]�������c|��vI�~<c����֟	�<�k���>�$��S�|�~�6s ��нD��H��m亚�x�;�Zy)��f*�S#��,��a\��`*�cxs��ƪDD�u1���=����/��(��3"����(��3��x�3ɻB|Mκ�
�Ӊ�9o����>���	1D$�OO�@�@1.m�6�A��׶�W�(�0U��#S�?Or"�}���Q���_A0ɂ֠|����*Ε���-�k���@E���	��{|����g�8�cR;�.�B��O�/����m%��pLxODGL�4����r6ؽ*�5�D(�ΛT�����#!��,^|F����/��� ��eT�5�~�u�Jv�׮��~C� ���y���a���X!2O&y�������- F\o��E�wi��B-��Y���#C� c��M�Js�.Ǖ�ġrɏ�H'`��ʀ/�p~h��<W{���E�R�o��ߨh��1N�Z��j� Î��[�M� �֩@n����6�����x�x���֗��Q֊��J����Ϛ����̼�p�.�? 4�'��Хh�L)�^��jk �-�e1xX�A�uk�R ����7y��D��_�j#D���0��y�˳�7��4�R|2B�ڒ��Z�����O��a�˶��1�|i,~����I��A.�ǉ��-��+�d�io��샫?�\�OC���e�`�H�2�4_�J��c
����Y�^��l){�Y;���;�st/&ĺ�5�3Ҟz�ae���P΢�-�-Ѝ�s���!�Xh�W�l;~+TYI�#v�f]g�:{�`a�u=������=W���sf-�X�5d{�\��=kn�'[�n��&�����mg��6<���a�49�y%:E�R�ب}�btЍ�\6=j�����\�]�ȷ��}��UN���Z���ULC�[��{�yL�톸����9�9�1����-���T���l�5�+S>�;�<�ౌ�\.�s͙��W������Ri����{� �7�r�w�)�� ����Ne� "08�i�)�����'�R�<�-K
�h8 ��eF�rS�K��I��H	b���|bUGM~�P��X�
	*�S٘�=ܕ'+��<X�c��V�(�#��k��TRd'<�4�mꏟxJBF��X�0�J���.y� ����e-̱W'���t��y|�������>��|�xrc���ŷ���(�[�ɦ����2�c��ʹ1n��s
��U6��[X���~}���G�p�����:Yα�cW�h<k�����T���9ЂO�{l�d�*�����A9�:H��G�pI\(����l��{U#���mo����~P��ծ$_�8~F�>�dҁ�*���l�9�F��Ne��U�A"�K��!3ӥ:mz�S-�,*��և;�������cψ/M�C�p���K}��q_�OK|K����e�]�,1��̏�ok�����#�����&av8r�;� ���;t�k��g����w'���p�9e1�!-tH��}�nz(#t�V�kܒ[Ћ�t�����jȄ���ȉ�ډ(7����b`1�S�b�l������ �eU%l� ���X��o��S�jbqlZ���W����:�@
�[�4��}{w+�J��QA�d�JO��a[��/����r�n�5ՙ�����rWs�7B�h�1x������������A��<�|�laa�f���FȲ�����^d���K�ﶩ(����\��>�IՁ�JG?(u�Y��yj'+E��bm[�E�x�!mb73B]�3�ᷭ�������}:�~W,���YP2�D�?�:TSZ����]F�I����[ƍf��¡I6�2@��ޘ�(x����.
�=�Z3z��0�3���.'��X��fSO���&�G(�&�M,���FK�d(?v�¯�UH��Կ�u]̲ש�%"�/���ڹ�#��S_��l��J��t0�}��`�ɥ���(��f��ʨ���@M�CΚj�R� V�'��Őd�~3�臺�*��)�sL���I�|��O6��!$�҇�Co��O�>���IR�z%�n&B����
� Χ�^*���f�.�Q���r4�q���y��
"��D��[\��8�	�0�1��C/:�ݦ]���M�D#/��-�
���� o�N�����_ZV�Φx�-UO�M�	�T�M�#w��c�Q䤡$/jʪ$�y�2,!����	C�W*_� ,p��:��A�͍T�Cr�OE��(��tF���8d������R�@���1�ѬU[T��|Xm�rR����L���Y {��3��P�g������u��Ӫpt��Bk+��7�N0��w/Ւ�]��.����{�Bp3�0f��L������)e�A�5���h�{�sڮ��ռ�.���XJ�l��h�����#s�$�^ܨoLu={ n�"�8c��ǫ��߫!�!<�<n�4�v�A�l{��f��c��s<"�9��eO�u�/D7��e`Zf���Bc�~��c�`���I�7r�H�!���-��V�YCW�9MƊ�.���Ld
I%�_��U�!m�lv���z�@���<�Ɨm��42����JQ���)��D�Xay�����H�$,w���sCz��Q�CVM�H��Q����T�^M����F�F?V���ah{��d�g����WPU]O5�93��2鞰&n4�a����|�}�9�_*C>hIU��r��zw���շmG�鲈���m�Z5�rY����'�q�|d�T����ɢ�1s\Q	lw�iGI��Kw�"(���ܲ�X&�
��'�I�ͧU�p�0��>�0X��K��d�
�-쪕���N�i��;�T	{b�3u?>L�J�Ҫ�e�b�O|UFp}���a������	��+Ԅiv�M@z
���u,v�=���"/�];,����1�jy�i��-���a��A�_cC�n�8ƍ�vr?q��y�e_y���E<��@��y����:��7���r2���&�]���9\d#�]ZJ�>r~L=��j��^�?ޓo�2����l2z~˴�����gd-U�ٰ^�������&�(ot�ò%q� ��?������c�0Z]����'�?���\��p�,��rUM��C�I�k�^��ϪN/���j�ݢ<E�\;czz��[��FV�3p�e�*Г����յ����)��m��H�{�!�H��8$p��=nf�R+���R�fg�>O�ZVt��R���8�ٶ��mUG���v���P���|fS���8<�H) a�n,����Erж����g�jZ!r��qEu?o?c%T4�i�Q �)�����%�Ճ��-�x�!w���#kٟ��ZX��Xֱ�c���d>�����tw ��9�-���fw-B9E|�����P�����ܟel�[�u��P?������sˡv˚�茞�+vu
�-]J��SD��=H�$�{�CKOʤ��2�(�;ȹ��q)5b�x{�_�cw�]����:�'�!�c �y�4�Z��T�߲�⻴H(����塆ņ5����R9Q7Ge-=OumT��+[���J�I����*q�|=�==P�+�L�$l=�.������2����d4L�-ĕ�9?6�6�^4!@�<��[�t�̿eI�`���%���PpIӨm8\����RB���T�N��S���x�@��s�
�<���"���^K�����o�:Se�r����Z�+_Hb�����c�����sJT���`��E��&v�oӢ�������TH��JYzq��RJ�3�/�>�y���f��yyYJL?�����B$kt?]" Kcފ[
�"�)Z��v?Ć��-��N�I�Tx�o�,J�w�J�n�(�8�u��S{�f��iصf������4@{Е2�'s-�fɍ�����l��Í�����RS� ۂT�����B#<���9n�I��{�������F���#ŚiG�?^δ����K���C
ܰ�����Zh�j�o�M�
����S2v�V���V+n�X��a�e�ׯ��½�oi��uO����Q���`�׎!K1��!�}|_��]��̺����r�ʙ{����@���oU�dƊ�P������h�y�n�"��c�����kH�)ka��/Z\Gs�r5-��["4T�`��N�aլl䱀�tE;@`���ۚS����bp��[e�~��c	�|	[]��h ��5D��C��b����:��e�-,�տk��;ft�:^G�FCq�y��=tPK�������C�E�4�N��r�ZGi�[��&�m���Ѳ�s���7�,����@��de�?%���Y ���3��ˆw�؃{z����$��"<�$>$�i���*���M=u�Ox>Mp������ɜ��[��2�	u�,�3.;�>h����t-
>����ʬw��L���orVj�f����9�!%c�e���Q�?XOp�+��ؼ�;����z��ƯH>B�4�*)�蚶f�[W�j9t��A���l����c����t@�⿴肅c�g��$�zOJ�:��U��F@�a-�Xv�[�t�$Q�&R��c�M�	+s�U����w<�T�A�)�e��BR�u�kC��c���=����l4ת�x?V�Hb�k6*À�ؼ�w��q�|�$�P��ߎ�&�p�!T>�7&+!���;��$�BЅii�t묽�=��|��"��o���bB�wsP�J�:�u)�$���L�ݟ]� ����9g�a�΃��:�6
.3�	q���z��B��4�)��f�կ���S���s6�������.���H�^]7-F^����Q����Rcmx���GK�m4���h(��}���AT}���w9��k	a� �x�$�-��WĽ���r>�w:ή9���:c��.q�9xԐ8���B��O"C��V�J	u9M0L�ܐ��C>�
'��hכS"9@�U7�V���M6�)hxX�&���.7E*��=è�V�d{&M���. [�A�8���ף
��Q����:בQ�
Vs~\a��}Q	�n��4���7�V�+ @�� b_�����|D���� ��Rf�u��3� fl�+��c�B��?ǿ��x��$Gz�ں{��75��X�s�,!��I�'���ՔLr�+l�a������H��&0<���
$_���ca��[�T��i	#��>��ϙu|j����p�%�I�f��u֧=2��Re&�y�¨8f�c8���k��!��u��dFy�ޔ������YެG�\
�)���4z���Qe�+�k�-�2)W�2�:��{�}��(_�'�,�I[�ϵ75�]I:[�4YIx�c,�*�+�C�3$�ѪJs
�������2������دV+��A�ge�ߗ۱���� �*:?1r�����82�Ç�W�#�~<n�����G�w�S<d����TO��,�w(@�!�g}RC,��I�0[�'Q,r��Q�.�
��^xZ�.�W�M��1���̘�R�,M�$�!P���r#��6|�V�YW�[����=�m'�i��?��E��v�0*P��:�G�$QC����_E�
�Y�K$%}H6��US�u��;xBJ�����qի�T΂��6�m6�"�q�$k\߅�ֶy�8_��w�@�a'������ �!P}!���+��v�B�D�e{���D���o�,�z�GO9X�a?~�h�puY���1} u�y? �[���(�`�6>���g��Õ��R�f�Ϧ�4ɍs��,��IfG��
s�,zZH |��l�`���nNy���:��xySn�M(�y?D�ΰ0���r�z�]XYt�c�l���x��B ��֗�R�LC�@uI�1m���1�Ņz>��E�3լů�ec�Q��rѧ�j����pȫdh&*�������-����.7i�c���KۼS�����0��Ǽ�*�/vHK4|/+xޏ���O��4��>*��6���~���K�V�!%��q���jS3��-�呿/,X����4�m�^����^�"��cP�F��S�"@'X�<���N��r3��ߍ����/��R�O��9���.��W���`D���7�|�����F�˲�{����U��ck�Y�C.�?,�r-ItNa|_r�WS�E��qmX�0OΨ00���G�y����P[�	��U=�R�h�>��ً��
��F�tf��b��3�b˝�����ū��r�tD�9����J/�m�26���}���o��+��y5LTu��J�#D�W�Z���귰���`ooV��)�s�Iג.j(�Oz
�Ӗ6���sӴ�������A�𙴋c�J�PF�Έ'����O~Q�) lЁzy���U�F���m�|v��@�hU�e@#��P�t��D��T��"�	�ڳ��8�8⟨!s����q$��3X4��ø Q�͗����H-��5 h��'���<��{K��G`�)�a��V&����J�:ǦJN���=�'T�l�(��H�>�(���p(dAhf�b�ܶ�y�f�?�ZA`���K�65�f|�B7��g�ړ�$h{���sԖh�@�7��씒�}����q�m~�]l�R�}Ҧ����t��l�i}�s���q���1�� ���u����!7V�2P�O�$��4�`�ݿ�5�h�/	c==��j���S ���v��5�����OV�rDM���S6U��7�� �zߣ~>`ˑ���
�ϭ���j�6�L�N;&�CI�T�tYum5�:��Q�̕Y/MH.2}�Mp�P��s��=���a�#��!������?�i��)Y^�{VV=��)[�����T�0�>���()u��d6��7�W������~Qhǲ>�j:�� �}�r�g�浪��Q�*�K�7v\�U��9��5�����I]�/�?����N��d�RnMड~rc�QJ�6gHu P��p.Sj�*�6��C��%4;I����0��YZN=�~N��Z�_}2+Ô3�|F���"p���z�0?k�F�3�zi�-WPDz(��5Ň�E���0��;Gr��E
!�E�e��;��S.R��Ǖ�O9�KDQ#aQ+1ӊ�1��#�Ϻ�2�h,E������!qo�j�V�4���k������lnISޤ���Kq@n��%�D1�<�P;g��@D��֫9�5�J�i�O�ʷAO{ρ���c%��v�V��*�&�62F(sA
!�3�5��n`�xF�Y��HC��o46�&���]���A�O�6��r_��p����݄{(�(j�	o(��Vz�U. �oJ�g~��C����[�YBB�HD���	l�""X��}���PQ��U�f�"�D�RG��Fg�;&��*������_��tϋ�P��k�	�v�ӐJG���Pl�{>��T�������ڙ�ݓh�MrH��_�w�u����\o%�M�~v� ��]��F9���vJ��[+1d�u�-�/녛��8����8�l��Ŷ
i��Y��u=S��8�1Z-�$83�{e%:����1���9�'��c1�#QH��,	2Q��LHܒqש)bM�Pgx�F��9�y�7�3�Ð���ޗe�|��W���;/S9oP���������i~�xtN�kj�۟oa"5z���1����O�z#�	�M���_ߨ�@� KVb&�~7;a����y����-2��u��Q�9O饮��Cwߋ��R����O��W�7j&�o|��/�I݋�kU��6��[��Z9�w?�5*���dad�f��?�0�D886'j����B��B���h�j�өXX��6[|e�wY��_�Z��4�6Do�_{TK�����G�iGT���QA_2k̝�,E����R6�~P�&�����Xee�;1 f��'�_���-9�ut���e7m��h}}�de�n3
�g��|�|�2�|z�j'�k�WIt[�����t��B
��U�Ŷ"➧Y��h�^_x�|��CGH�zl\-���3Es�X��;J�� d��4�Y+��[{�
�;�����yzTs�>������;�R���G-S!�x��F���O�s��Vb�h���}{5�k�]Wo+e'�Q��bߚ�t�[��l�����l�9u�?6�S�|�����f���B��YIF�!�C= uz��PĮ�R���g4�<O�|�Zγw�J\�<�ql�{�ڨBNl,��Kp�X���HF�q��Q��cW7�;����ﰵ����D3;�����93�qG�z|h�8����{T��6�|^u��&n�[�ï�����v�l�?+����P� _}����.�2�����њ��/���p|q=����D��.�S���i.\���Ya��pN r����t�?�($�Mb, ��@>1��^�/�ڤU4�[t�|��JL�ߌX>��I���ݷ�1���c�CB�Q�;����}7��S�������jPE����{�Oܸ�%���\�Ç��S��r�[��nے�e����+���9\e(��o�d��*y,E��V�O�Q����I�nL����w�d��i���#o� ��I ���as��,ę��+�g���w
�{²+Yj�(K]U:ͷ�#��>./�ɡ:j
��鲎�|iMW��)���������u�m.���U�+⵴<�S�<hJ��[��v.+�#��XT��kI�bw=O25����� M��L)�'Θ�N�u�w����Dd���Z~��wd-\�Pd5� ����:�TP����9�V��������εh)Zٌu��jx���PJB�-�����b�çL�����م��N��M��Z\ӝ�ef4�,�4x�wz^1��z���!��ح���d�Xl�*��KBH�a<�b:��Mz�`�%�+�09l6��EDd�=��؞2��S��l+�r�|�ZÚI�ef�2��б�[����j�:w�>�}>��x�<���K�@�{�az�0�-�#���L�ݺC��+��9�xD�s4��)�ދ ��~���v"�͖��(Q���	m3gBK�%�
�ū�C;�O:1�8Н�,�H��k�[f�'�Ӝ���B�d���~�$�6�ڶ�t�A
�ړ`���J���Yٶ��7=�r�4���-���j/��oٗ���Ki/��N_cbf"�f�Y�Ij�]�N�Q(�E��ZS�u���!%���V�t�ʼ
��_#��/
='�>��7q1�5S������o��,׻�!�7�H�U\T�߈���%��m�ɇٍK|+؋����"���^w`+�FA�u���&ف�_�8���2����!n�c)Cҍj�w	��U�����Xݾ%a0�æ8�EY�1i~�i_���แͯ����CJ^!	�2���L�>䖼?6beảR�̯NL�5�ƣ�Wb��O����w0Gj� ��u�E,�������+4��[5#�웂�Ȫ�bL*7ՑU�������~D��F���������/v�	�>|LX��˫B�3s#�.'��k�M�;��>�lZ�\�Q��t~��۷�%��@�Jݵ��"��Ev�"͎�����t[ ��k�K����8D.؜�ء�(#�����QC�`�����'ݩ���ȩ�B��AD�l�����L�/=����̩���i�T���]����?�T"����)��	j�<�ux�2���(ml,K5BQ�tҠZ�ɫ{���er��@�qYc��z���Z�.9.�J���	�ʘ��2oqHR���ph��ҥl-����@���.��񿲥�rӘ��
n�`���h���<���)g�㼓��8�c&ר�p2c���{MV`}9D�1�`��_kТ��;�@zG/��'g�ZP�����n�C�0�M��-��V��M����?ԫ�úw`܃\J��B��p#<3 ��;L�b�� )uV�7������������������X����.��:���Jq�8���$5U��P���U��,7�r��CjP\ܐ�Q����,�Q�\ܒ��;���U�?\P/�4�P��(n��S�Opo�����v�9���|d*���Ŕ��B�9� �������xǚ��k>2�hV��q�0߂� � /�������۝>bX�3�=��'���hl�5�0�Ϗ��*�ŔE��c��G�8�v�Q��iAn]�zx��J)�]b�J�:J}t�8�����-%�L"%tս!�*�Ps�xR�K�7�)�i^�&��D��D��̏O���b�O�X1�n>~�^�w�=� P α��x8�9���7֨$�(&>���T��	x*�A���nli��j��c�s�v���]���4E���o�� l�W��Y����vyt����Cs?E�OA[�?7��S�o��I��*��K:��M�S-��Ǯb^3��z��Q�kU��:G���mP!fH]��o�+mM�#�sn��A� 3hy6R��'C�ת��A�� zD���&Qy)�wv2/oA��dꭤ�rj8A	Ī'tR혍�Z4Sq���è�o-��=�WQ�}��'w��g�/]��!�]ٰs�8̛��ak{��2\�ؔA�AQE��-%�񯔥y��y�R��k�LV�"�����X� �y݆X\Asߵ)���ر��Z�5�/�mZ{�C��\7z�V<���~�4�3��$�$���fUc�A|t��2�#�}��Dm���m����-oؓ�� >`��RR�_5�G�<��!��8�'��2]z^�xG��y�sF��7��:���w�w��֐;���/�@�Sg��f�����I�MHO�|�־eW�(������~��1/�"l��.�c�nS8
O4G�9QMxx�LR��kQ�&��p�Sq����@I;/�q#I�K���E^�NQ�bI��>֑��[E��9.i1���r�Y����ĹI���C��B�,�� q�pA�mI �;�XZ�Jx>�8����)��
���o�"���-\1$����V�C�����sy0
sK�Q
Ācu�"ZQn�m[X��@k�]g��I��-
�Zɒ�yxW�$����O��>Ot�����g�|�Dw�Z��AJa��e��8�ѼXv��[;0ӃG�d�/��loy�ʕ�@��zʪR�a�f~��s���>�{sV4F�wΗ³b�
����_?�3(]���'�W��p����R�H���rc��ME\� �F�eC�Z/�e�$��N{c�7�K�4��"�i�kj���c��{�M#�[�2D�S�CJ�g�0�Y
AGɸ�-3û�N�w�#Ғ!��V���I¿v=�D�]5쐮����=}uDғ�~�]v6�H,fޝ��[��G�o*����զ�"��S�n}��� 91ۆ�B��3c$��U�-ab/![r�~�n���g��IB����lsf穳�+'չ���c�[��	��\���:��,.=F�
�?��90p�?EaJx��ɬ�2�Q&?�'��"�ӎ��������9�f�|4lw��8e�����7mf�5��:OC!��+g��e��wߥ��5q�ͯg���z��r�|���v�����	ʰ����4��-�ɳ���߂��װ�F�[�"���p9*����4&
>�	 =�E��RظSC1��Qe�]�r<D�.��F�n��,7�x�z�!���4o�0n�4O���F�XT7��ͣ�Al�fF0��8^�P��-�'��SI:/%����Zq�R2 ��v	��#WG���	��^~��졘|X}_f�d�k'MdR����o��ʑrڡmQ��g�E�������� g�[ZIa��9t'�V.�QQDV[�[���|;S��1 Chh��T�0��&��^<0�ܪp�_�6�/��� Wu�(s��aN�!�Q��ö�~s�4���
j�Dv�{�=��ho�@�fZ�<m.zrx��z<5f0�R�1�A���`\�F ��J}m��/�B��cᥠ8�q�P U�C]D���෽�0B!$�e%3���F�/t�[�[/[Z�n�tNn��~�����ܝ��	��#M��� �RH�ᰏ�����dS�����\�h��X����7�աУ@�mڰ�gMa��fu��	Os�7�j�[b�g��\���#6}���t���i�y�g�߃5��2(!��DAxb��ʩ���Ϛmw�=7�'�������Z{쓽�=r��� P�엽�r�X�Am��:��.a��F�y|Ŗj��;�̺r��a��/� �R_���n�v�S���@|S"UO�ϰ����9{EX�� h���q�B�c�6�@�0`��h�"S�9������y'�=V�z�^�Nykf��tg�ТT�Ft?�����O��`�]�ߺw��4��;ެt��SN��87���2��KZ	O��Pߓ�O�Ё?�x&��(�t3�I��Hgc�O��W�}��u(�4V�;�{B�)H/fĪ,%�i~��7�^h\iR�M��.�DfԔ�K�HΏT������qs8�?��wˊ���b�ǖ$2@!�� >hxI" ������駗yƇ��1�����*=��)�Z#���>��yc���(:)�ǧn�z��f�GN� ������OX��P6��c���+��/R��\Q8J�t\o9 �L5]1ø�	S�R���v��`؄%'�<�Q��8ń����A���W�^@ǲ8K&m�2 �_C�R7���-����zY2|���7��>��Z5�+�0캾A�!���PcKpA`��X�<��'�O��YI@n)�Pi���h���~����Ǵ�J�p���pt���"����d[j	 ߖ%���BSM	��O<D�>b>	RB$�}��ـܙ�.���G�m����� ���R0��d�&�Z�ي+�/���&K��"����V��λ����t��T�
�s��U'&�ye��e�T�AK�����(魼�2+��aT�?#j��q*��c���D���gK�=�8��/�!�Uչͣ�_���zB('2�K{s�U)m��\
�Df��z��d0��D����=��.��R�i��H^�o�����[^3p���b��F[}��y��cRا�K��I��Ko��c��	odl>c#��� �H��J	c;�1�ت���	* T�C2�kz+j��ɩ<=JݔA�����O���y�?�֘3蠕w�+�O�0����7w�^�w���οa�I�6����C��O\�,���&J�ɀ�-��,A(�|��r�����k$��N�*�G��Ȩְ�t��f�8�ӯam�xo�@���F��R �Z/	�����v�se{/+ओͤ
���JՙUط���,����fc]��%�_ƿ�:��1""'��Ҧ��A�J��w���z��.����A��S�f.��@u?���^������C\�7t۟ԝu꣱��i�^���l��Hz��S�)89e�Y�������rz��F��O�\��0Q�y�tkE��QX(��w����{9/b�פ5\.�R�4i��e�zH-AWrϫ�iN�[�нPW�C�(y��xpLEW�X�� �¤+i��0o��.~S�[m�k{��ydJr������'Ur��+-Ce!�}���5 �����I�S��� .F?8}�ܡ�c��9�B��E󤈇�P�A��l 
�M����J�JT`�"à�d��;K�<��^�Z	5����,�@XI�z-���VqNO I��I*�Ef�e,���38 Y�$'�C��>_7R�7��i�r8SpDv����5�uОC�K����p�穁����_[)|��i/��1^�ץ�?��3J�M�3��]����\M�8R���r���	���je貰�B�ϓ��L�s�ɀ�`��VA��u�>a�ᵜ�e�@��0�:���΄e��iɱ^/���Al�Z��>Ӗ7_��}�n�.�T��h�K7:��F�c!M[WGc
�c�1�'�뾀�C��'E�lƳ"��&#]�������7a��7s0_��C�ҽ��R������Y�98��U<vr��G���y������i��Q�X�K�3��WG�����S��X[�׏�ll��&ڒ4���m��B��]��tr�S{E���/��_%���b�H.���e�zwY�훁;_M9����7\�#e^��5�����zU]����j���ix�}}��M@#��Q��K�op��&�^#|��T�k�� sh0�A�Q���)�	�-�ӈ3��s'?_��û[Mʹ���q ��w`�2�d�$�~$_�*��Z�t��ٻjk0�z9Z�#Z�XF[��m�!���ڃ;����Y�9%cV��k����գ�+� {+�وY*.HD��8r�+�ޣ&�s�����m��AרԜ��bkן��%���W������d��W���I~ǥ��V�Jl3d����wf����.gxAڣ��{���ϻ��S2_��9��BFѭX�:/(��!����^��"
]X#]"�I������+�}"k� �'~x@*"D3G;2S�#(��+��snR_�KzQ���{��X��m�~#������5�I*��!���`CA?�(Y���/v�I�u����^���k����K��������r}ܠ�-2���Ņ��m��s��I����N�$Z��MD�4�Ds���A�J�k�B0O��y4�]1�=�++=��|�C��z���Y�F�Vz�#� ������4�	�2j�*�l.W��Xw��Lu����t�;��``ko*�M/X	�3���f�b[�g#��^��b
���K,�J#��Z�+�����4�1�,У���گ~������`_eq��"Y�9�Q�֑S�΅��A���^�i7Q�c�F3~�[�+db�� ]�3��~W����_�S-H|�L�^�������mJ��[@�p�T,|��S
��l;�+r.�m����M���I���ˡ��LR�lg��:�A�ml�S(No, �$��dD���ݐL���AF
��ث��u�F	���������۹�r�#~e��2�	G�h����h�w��q�\�HwP�Y0��3��K�{*oX�	iՈ
&ɧL��|���&	��%5}�9�/���xN����ܵ��E����yzu'$�@Vb��}:���tz��6�"��%�z�%��)����{�����x �e���d˕^Q��;�3��xm�-]�Gԯ�h�Ni��
�0��ľ2�lA�������*�4e�����k>��E�*cw)l��댪��
��y�G��y�j��VI�1G�c��:h!�Y��H
bf &�$ٕ�W�^�_)�A�ze� ܜ���UӍV�'����x���+5�O&hUY�!.d/�gh�H��V�V/[�(��r��lr���4
z���">�Z}<�Eup4���7ʢ���,��l{AYp+E7�D�_g��I��C3GR& ��+�;�����pOߤ��9@lp>��ڧ��0�y�b��?���a��))m���"�iS�~��5=�á�G����rEcUu��G���`�e�&�U�"���U�Ậ�{)�`���P@��b�)L�z����y�b�f|ړ"�X랏�336��sA��Afͺ�zꢅ����˴��%z�Ȫw�ƕ5�������c�V�'jj[xv�^��H;.;��W�L���i�%Ƥ@y�0�(P~4�޿0�x��`{��f����������^�]����1|�%��*,[5�|���_��@b{��$[Y�f�o��g�T��#ɍ�Š�w*?Fm�*��wI2v]��������)�`����i5�OB��h_]1\��������,1���6]�
����;U�s�ț���-��*\��� �*�G�n��&zv	�FS� {��N\ybd�ιK�[����.�� �ˊ.j5A�)"��|���3��� @|�Q�`�6�RLz)�������b�һU��[�N5�Mj~ �Q����%j�}`��%��&6>��7C�×���}���B���q�kȴ�CC7t`�D|���.O�J��`�=aݟ8��>��[�կ�1L�K����m�(��h#�:\I�;33�1k��W���w�}��xt�Uf��� No�O��%g��h�~���T9抆��ٌ��y�t����!n{��"����x-���Jc��o3�B����ׅ۽Vi{�n������		r�{�Y"w<�O�
�.6����~cq��j:�z���h.aQ}�1�TT�0F^e�����#�ǉ ���U��d<��G��Y>_��5}��7��t#S���:���D��n�{���.	ߎ�)!�����}����_O!H����@��˪:�¯'Sc���	.uD�U0
&��A�8?��|H��*��i����ޔZ�vh�-�3@�I�b��d���U�ßD��g��R;���B_,�2s�!��Y�Ɣ9!�؟�}�6JP���TgJjg�G3b��ĽH�o�\*Op9��yޘ)k�i�:jH���X�\^v'�OgQ4��0�-��
����_�POe��@��̨�u ��r��X�Fe̗�Fn�hSA�X�[8�+�X�"�Kr�$�P&b @�e�(*��O_�����3�DХ�(�{c�~QY-��l��dR��X��������?�<x+�����D�μ_�rt�x׶D�O�K�����,�& ͂��V�B��c{�[[LCȵ"�Ns��g�����$�]A�YV��Xg�t�m-��W���dVbe�G�蹜0��^ز6��#�Z�X����3��w�9���b��e4
�f�"a-}�o!+O�X)�I����/TM�&M��Y+~�8@�o�b�#k�K(�`B��rDG�JH�:Y�-=+#O��y�j\\��4�Qά/Ζ�HbJ3N~�N'���ITj0��*�n��C1��it��w<����h�|�]�p x������N��A�ۖ��fЇb\
�Ţ���Ĥ]D�L"sQ��� ��r7�ɗ�s<��#O�"��
��HdW��q�R�P� �٩b�ٵ�N`�J|[�v	"5��cݓba6i�"Ԟ����F�Ƴuy��ޑ �UيH�]4�0$&n�&����-XN�P
��kAe��֒�������Hb��`{�=R����g�7p�~���R��&���Lg�I#��!�D8o/��U&(Fd����C�f����J��cg����M�����}������I��s�SCq��o��7��+%\�?�A�PQ��es҅���x�A�7#��H�v��\�ҍ��"�F5>�-�����Aɫ�����NGUX�Zy1�6-߸-�{�Е>.7���o�?��\>�K
S�!s&�w�%ƨ&>x��]#��'>�0@3&�Ar/�Os���j*z���D5��[�:�=�]7�����~�R��h�;�h/^�E�z'+���e��},��f�qP ������E��!<�*�GpD�1g��d ������Ch;��c��ԶU�?Wg��O�R_l�ŉ�_ZmI��´���H4��%ߪ4d�Ua��(S4�A5��)�y�s�\���S<�7&x8�2���8����wk���iE��hU.i�|Sg���"<�P\��bd����$�c6/,Gk��N�����QGY�1ŉ�Nå[�T=GU3i�X{�����o��4%<I>:�5k��?�A��u����3�y!堄9x\;cf����d�������\��WNhN>�\���m�>:z��Hf�lQa��H��r�3�vv<�G3�X����;c����O�Ŏ�k_�B��^��z@�$ß�KZ�X�_d��.`�	����.fW)y9�� P���k����8�xyʃi�_\mJ��&����(��_{��-�dߚ=���<�����yE����'��[t\)�����i�զ��h����Ԇ��>Mj�s�"�gq�Y��a^��#�Gs�A�ܼes��KY�vlsq�^Ϛh��pį���o���r�w;�����'-����ײ|�97���l��`yӁ"�u3B�4��
p��R)�Sз����4x_���
8̳�f��^)����(YK�"�܇푷�QP�_�4�V7��蜞�5��v.Nh�;5�²���	I�q���?����&Ag]K������T�:�������ߟh�Q�	'~45�r	��zG�S��w��F`�z�}¯JU��	��6�aL��^H}�ѫ�����`y�i�;�I��Yi�Nb
.�w��ܵh�l@c&P񓙺}�f��*]�s�k��z����bݢ�1w%>=��o:U�\�� ��:�s5Q�7w�!��9-��G�����2�/{#�<QTD-����!��d�Re?��-G�Liy��5��A�?X�/U�[��D���}=����q��Y�5E`C�˨���0��<�*���[�3�Ik��:HÎ�M�8�|�">e3,�� ��".*Ƞ-+���2����������Ն�gOY^ZK�%'�8�%���W����sM2�/h�����ZC	f:�=��W�� �@1T�JS�*P7�}6}Ct��Wی0d����W�?��D'D'�6};( �yTC�͑�u�S��O�+�v��>�~���������c��З����&�{�r��F&��j�=b����\�E����d��i̡R�5��݆���Ya.� ����vqP�Q�wȢ|h	��^eMO��i���f4X�Ǿ�"bO�f@M�$%5`{��~�o�~��W�N4�����@�zn�GÛ´�q��&Y&e��௚\�������^ɼC:D���c��?���_��ۓ��&�3`��͙�t��8�9y�#>:� �ق�$�
 ��zSI�m�![�YT��3��C2!~@�={V;�=򮵕X���^��k�:�sn��������Zn焼��)7��XرH�˥�^�W'��)��$���+�A��ZA��;�����-�.�w���f�5-1��PX]c��.�g �2��+���:�f��r��fNW���ba�Hd-���X���Q|���4p�=vs
��q�$��X��>*�w���H wH��.�u�.�^���NnN�$B���gd"JQPF]D3�rjR7/=�C���e�Q�"g��}�,z��=�u�C�����o��2<�䚿_��βLnO��aq�a���!k�]h���Z����vm�w��n|���F�1[��+��ow�D|y�;�����c���߁h�b�ʔ�.���9��h+�X��ϫ�o����J�5�B�KJu@4��%�(�/�*(ͥ�X�ܠ��m����d�杉Z�2�b����m*��O�3F�熀��HasC�_�����Ն��}n���u�1O�-��
]�����Y&p�ӝ���{3�yGt�d�:2�M�����n�PO0i'.N7?��	�ky��鄩��o�l-
Y�u�z��P6�V��Jq�
��A�Gܒq���L��]0QK��!_
\��W%r�e�k6�t9��N����H~�N]�"�c_����:Z�������`�=�)���X�z�3.�N����-���pꅩ[2��� 9��Yw��)��v�����6�4�ӭ'��+�	̠�Jo��s�x���|D�z ]���o�?��M<�}��l�H�*��(q)odv0����X�z� @�⃏O�Hc� i�C���!�W�<�< �
C9(��a^q�žʼ�?���t�j=�f�ʪtn0*U\f��f~���|r�
Ɲʋ����::
���@�g��i>�ɲ�(vT/��'J�$�%�7w��G&��I}������:A��)-A8���=�<�љ[FV��Ck	��LHn��Z4Մ�Z����H�&���V 'y�����ݷn}O7���v�Z���9-��&�7���qⶳ�U�h>��K��t.��,@g�Յ�(�����{��i�Jp�d�,È?)��,H\�]!xO�#=W� ��g�L�G��D[�Wn@�����������5TJ��q;���ՇH$
��^�%ѶonYu,K��&�`���B$���M]��J�N.�K�7*�J
��=q7���먽��@����{ ��'+	M�j�U"�#F��c5IT�&�<�H�
�KԸMhR���O�Z�WFb6���,Tf�s|ˡ[|����5�|Ӳ�%,�a�N&t�HOR�b�~��C-M���d��h�:�_�>A5Dy�^�fJ�Gm|P��q�`xEh�s�=mw(W����<��sL���Hrnn*Ń{��ղl#ue�!��1����%��n�{ax���˴כ��)��-i��e�%F!~���E=����p�PI/}_l[�6�Z3�I�)½�����%❕2���_.'b����)���V�Q�_ЪbH����4DJ�`��)���bv.�i�F��Dh���'��T�������8\�=fY�m�V5�i�C\��N����n��"��� ��<y���a̤�-ʾ�'xc^��n�yrW�?e\-f��b44il#A~�XQ�;�MVc���w�F1v��J����$(e�Y�p:z.2~,��M�P�UG��qb�����d�鵁Y��j�AS��c,��IYCu����P��y�:�#���Lt��(@�U�|ggy�a����kǕ��]���L떌�`xcx?����n���$�1�žR����p���5�,�ECgSP��x㸍�&('Ԃ�b�L[��F�q�ɳA�-��a�HW����LWx#'���E+�H���W�,�;N�Ǉ�"�!p�4�Č�:����'�����灐#>�ݝ���n+x�3���>}'b���� �����q�`���~xT�CQ1���h����~��c
�h����`ht�@�����P6D}wr,�f��f޳uo!��ݟ�DY�`v�V�<���>�j��3,��u>��C���U��Z$9nbw��u��(�U�����`_���*#E��P.�}��{�@�6_�w���9k��R姀Tj��v��i�GR	K�F�o��#��t;���Aܦu.`�zGi�i�tX��t����v�R!�B���Z��l��K���Y�td�t��#pcb(�i�<�sʌ~%t4�Ŧ�gC+�+X�٨�)[
�j��9���Dfȯ�R��()��X!�$�����L���D�)��<��\��T��z\�3UR�Xr�Nw�Gc��3�']�V�)FҌ`x�(�&��f��Ϯ�g ��,a�X���P��:��"�٘&��s��2���W��9�&��d��p���q���R���(��3��9��=�ht���}��H���'�X�Y3���[3T��k%����l>)hOs�er��Wi���&1I�!��O����������[����l�La�M0z������m�rG�t�8���:5_���2��[k.����x��^���E#V�G�8v�vg��8��+H����]�4�iKΎ�0�dl�讈2�pq��ɯ�.��z=!>~�|�K�;T/c{�����L+���/�w�:86��\�`�'�3r�@�ƘP|�ҿ-��7�/��x�L`�?���U�S/R���=@R)�#�2RD� ����N���b���fU�T��b�^��������B���g��9l=���k�r��i$�"��6~~����e{9i��%<)��|~�U�C�d��s9>U?^K�Z��pm�����PNAI�����9e�Vټmq�9��ˤ���uvU���+b�&�0�������6n� 	�����M{�K�\A���|C�CnƁ�)��iϲ�n�cb�(��`���Z)��z��*$鋿�𞜂�{�����uV�P�ܘ��.{�+����4����PVQ���P�2K;�s��?m�R]�H�C�x2�y���4K�լ��zw;v29f}��o�� �sP%��ѥ�@��<��;�!}>TAI+T4�DW�`���;��Ώ>܂�L	c�M��A����aKCs����+,�M�I��/�B0��i��/Ŷf"����7�>�L���$
#g^ذw��]L��7���8"B���+��hT��ym}{���p�
g�?,X�aJ��=�����!�����:�;,/��א�j�Kz$�F
�E��a�ؓ;%��]"�|fQ#�|���u�CA�W9cU��Y.�����U�$`��{�'8�I��<�����~�%O
��X�w�V��S��r@�]?'�~Ō�v���i�����y�6�������
?�f��4$��ĕ��ܢh����.�2L��id��Ҡ/p
��E����Z{3���q1�������ɬ��͝��3%�1QN�߆v���>k���:�XGh�a�n ���"BD�#
�76�陇�����Ŋ��n2��^}�]�����gB��
��7��L��@|1y1�O��q��(\G8м5��`V��]��2���_u����f`�D��.XC%�P��F��>}�(�,ĤS(Z{�ظ�� D�[��m�Bt^��������l�Y�	����u��n��&RG�bT���-k�0C'@�?�X�W�`�?�qD�|�@��E ���{�)�`�UΉ2��^�mA�=�|��Z����p�#r�}����z#�/Pvk�����M���eQ���
�f���W��UĠ�H�"��U<�Dɝa��c�(Ϲ�(�o%���l���.��
�������]}.�L�O���*����K����W�k.�iC�U���:],�i�}��{N<�	.�Z0n�� �K3 �Pp���>�d����i�
�|:��N[�s,��a-�Ű��O���fd��pL�j�����4Ťx�q�(��~�V!,��D�w�]�+����$?u��܈�o���aq �-�B�-tzo��<�4sJ����R��q���Z/ƍ'�u��x�W(_�n�찑tRS;�ߕDLP��W�z��(��38����^�vb:��e��a�d~׏�s��X���fR�Ú��#�\�! �^\�]�CY�z�q7�V�g���6b�0F+:Jbp4B�S���y��F%�ڗ�N�����/�X��z~< ��֒K0�s��}Q��}����FU5��RƎ� ':����g�T�+߶F�fϚ�o�oӁ�{�K�2j-A�����)6|��[���꘬�u>%���q~�$U�6D�E�`��n�.v�	?�;0���?�nZ2R1y��+>�����-�8K&z�N�L�e�P�y�N4��/f�j��>p���L��uo���坥�\:����)�����+Rw'y]ݨ?��?
.K"�GKe��
o(�b�3��ѓ�A�<��xi4�S�{�Ai�����T̃[�Ќ
_J���j�+��"v�����c���LL`n���M'<C�U�o�;���#[ð ���y��l#�:�l�Nk�ߒ�9:
G_b���������	��s�`u�%�����7K���/n^\gH%��2���OV�(7b��:��&n��22����3����#�>I(c����ר�2#�xE�Х^���q��$�/ݤ��,�{8W�KT@@�-K{��ԋ���)� �f�^�2�pۀ(�M����f�Y�B�M� qάtN�ч-�3L��6Âٴ)���W	1�����è�~*ǘR�[��UGo�t<�~��HC�8J.ܮ��4A�9�^�ֶ�I� 4ؓS,-Q�噮O�{9����C>,���AY"p��%M2��؍/��zb�X�+H��uw��ac-sbCגT��4I��w= B6V�/y0<��_�HB�7�x��'v�**B!CBR��A�����tL|�s5C��a��z|m��7��ƙ�D�+w�<�e��L?dj������a���t�pם��y�E�,�/�>��l�������M"A�Eց��.�������
fVx���-�K�et>	k5���1g��L�4��8ੌ�g%�{�1���P߷�)�_ɧ�L�4a3Ȁ��f@M]�V�z	i����,�p��v������B��~�^Xc�ѣU`�BY�l_�K��1<GV��\���
��>8��#�^�����_�ڕ���w-��(�lz��i�J5��,�V6�L�-J=�O����)��Z��S�dFG��W���H�A6��l��rW��WjE�䀶�(OS�|+E }i"�P�-�����𨪇i�ψ�e�K�:���L�	�R��d���G������׭i�F±(��y3ۉ�;��w���[F�/�nɋ�A��T76��O�Ύ�Q��?������K1"�� �����!��ԁ63���АX9>B*�����Ł�Ls�vg�l��I/Zci��ոeE��d�x>NB�������
: ��.�BV����[�Qs �
�UFڝ�e8k[�rI��� ��c=}ⱱ���Y�0��(L������xR�}�š�b�������f�2�Y雳CH�h�ƶ�ˈ�4dG���\1�Q]�>�zZ��aC_"L&$=���o"��ORz�G���M�%c����3�8��;Sv ��n<����O�6���Gk����ퟓ�-'�7Kˬ��M�4K���3�2O�t"����%X76��m�0~����T�L�ʁ�F?�H���.�?���~��������S2�Z�n� �����R%M�"S���Nѵ�ۮ6�H������ ��Y����Z�(D�\G���Y�}I��ـ0ǒ9���kŪƄ����T@,�j"�m�*;�k�]�75T�Vo��ֱ�.J��OQ(�a��������*��VO�s�_5_���h��	��q8�5u�3�bS8�G��PY_)v��%����y�
O�a<�9�0�um��2n�>k�	�i�	���s�޿���S��EZFihs���Q�Ҝ����(���]�_<YQ�|�k�����O�쑹#p)PR����
��[9	��E廪gg��]"��s�
� H�@Jd�n���i6}B�l`7O��r����5���᝘�����I���~�r��J7��Q5x���jK���z�3x8���c�4�z�̫�)e�reO��@���8m��|Eb�v�!�Ɏ����]}ꈤ:wT�mGk�9���Q�id��3I�O�Q|݊�	�*����I��=A,`��Q����_g�T�I7<����)M5a�J+��E��~�:������R����)�� V�۹.�\� �saq���A���*v~����/i�:170r���
�jh$`���E3rus�	�Y
�9��%��a���M�Y�ָ�Z�/O\Yb<`L�dq*� uS�g7pS>�7�mM�NW[�n��9��f�]կ#}K6���JH)�E��!A�F{64�^�E�{�3�e�x������s���7I�ަO���m�^v�kI]�J_NL�K-ȶ���8�A7��{�q����' ���q�&���K\W:�p�^/�$��7Vʐrs�^�Q�6yD��YHlN�MM��-@,ü���cnc��*~�-9v4æ�=��F�J��XMDH�נ%�wi�<tS����h��K�畝�R�D��Z��%�d_���4���)	�=%L��3{Z�އ7�����G��������qF[}�X.8n�*���l|.��i�����݊:.�{��J��m�*p�+�����@`�E�f��"ˊ�Օ��i��^��RZ��Γ�fZfݙ;�������q�KG,�Bl��v{&�K~⊒}�6n���J[̮�ѲU���֩QQh:p�Q`�^��)"E��n/�-1PO�-(�ct�=q7�S��>QQ� ��<t����������U���Z����:\ֲ�Oϒ��ٽ���[/<*��$�c����v��EC���.J� s�N�82��p\���o�CY��leM���k[p���Ƕn;3�D�m����O�k�R�hg�6�g�mvE&���\��ڣKr�l���k�
y$��"�Յ�*�� �t���;�K���8܅�(A�>�rsˎ����6��WGQ��L?���cR
'�nYǰ��y�ST���I���̐�Y2_�͙(�4�N�y̚Ҙ��N�P�7���\=
�&��Ӥ����_�Q���L�{���[��0P���OM��'�Vf�a�E�N.~��u�H�/!�����+�V�;�&��&����;�BՋ���U.������&�GY�.#�	'h2�U?�S)Nj3_\�"㬬�����Z[ľ�py��ԫ8q6T�ߓ:ļ�5�&%p�F��+L�?�&gL�E�E=�<Mdݔ���oy�n���h[k]� (���q��..o�K n0��v��2Tk�j�r^@�ռ:=c�K'���ψ�MS�i%�5ȼfx��J�<�@ 1_v)�1��ݜ�;�����@l���E6���rH��nњ��p�)B<el��}���� ����.�y��hcA�uc䟄4�!�歷S��&�U:1@��}ސ��ҩ�m�i�o+u�����֩Duq��5��8��8^T��<Ol���o� ��p���}H�WKϤ��$�B��W�¹��ٞ��kR���!���4�$�@h2���t)���T\ [���Zhl6�P�עԩ�8F^F'9�է9p���0�_u�}�Ѕ�~��F-�3LP�I�~��r���jI��r���!S�N��5�tZ�Ä!0�81�-E�ٵ�E$�t���)`�ܷ��s��wAV%.9c;�{w���mJcԙi��B+i�UA�����Ж���+sC�^~�SLp�E*Ӽ'i.��>�� m�����D��|l0F�=�r�;�?ă��~�/�W�m���r��C�
�=��#&]
D;��f�;I��%?�#ǻ�OҔ��� Fz<���W<Q[�T�-�/:��D�(khq�v�Ԃj��QN j�:Ч���x��^H��2��n�l�ò��ub�����2��.��ǆ�޸��ZVYCY���j8���\r)�	w�U��6:x�����cZ���@Q4SM�C[�U�ZʐP��e7�TA]�_�7�]�0:d��@�~J����u\��|�������J�fw��w��Z�� ���^5D��a�#��D-�1�'�=��"��'�I[�{j��e������w`�	;bW�{aVK��s��?�yd"@[����za��ڏ�����n�,�G�p��l�/�τ~"�<�H����7����:�ۑK�E��������-�1�+C��D�<���5����а�nm��L�����$�Yި
��"(����I�C��a���u'(2:Y��׭���Y+Wm��o���Ҁʛ=A�A���v��]"�,�h�d�n�ǜ&C��4����U�}A�v�X�n[ey��wl"4�ý�%um)I�,�Fj�G��!E��?E�%�ߧ[����?��BBe�	6}uB!�rv˃@����2��P����ƾ���1�����qo(��qdó�/�|�K� %;�G��	1iFl�h��f��q�.�Ua���V�� �U��" #�&B���YG�T?�d,����4��O˙m���8U�S�|����/��+
��2
�z��r��L�)�8@��ر% ��м��M�_2u���������b��u�C�j�1ͼ�J��p���
��s�	�X!F�3Xj�y`�O�.£�sX�W�R��fK�����D�e��C�p�џ;�(�p4�5q�7�?'����9~/"���^9&�)��'�Pσ� bt�Ҟl�f&G��
X�+i�����C!x��M�y��+�\��~L���i�~�{�����٦��������CeTo���(����6���e_�)���T��E�<�p���t`���6#v^t=�L/1�U�#b�~�Y��u4�}��2�% .w�VD�/�����ߪg���Z/�����7���S	��s���_�����ެ6��ի�K�z|�CPk�S�b�5p.m������S�����k*;�E�|7Q]t���#8=��6�Wй6���T�V~DbK3�ᐶ1C�?����hMSn��&I,U	���|�=�א3���!ڀ�'��}�&��ڛW���i���/K>J3 �Z��â�������'���<��+�E��4,jT�����{A��:�a�bQ�^���Q���"�|t�o> �i��� �&nbOm(\���S�3�7$�0��qv�2옩y�,��(3����Jz��n���,��Gn1�:0��b�T�LlR��:�u0�4-I.f�)�x5Ҽ�:�&�A���@��yQ�!*�8���TBf�ǜB�7��3!���{֧D'�Q׆A�m7Z�*��.���kO�qG�@�G-Ҭ!C*��Mq��| i�B�{�۠�+ �T�����Y���Y��J�gl�u���� ��A~z�d#�M^�	� �?���ۂ�A&���Y~��/���,�V�7jF�%�J��ϛ���|t��p5��~�X	��Tɴ�.QF����U�dD�5�Y%���]�R�.�pޏ8��jE~�I�uF-����G|��_0m�T���[�e!��&� E[�k_-hm �"2�آP�����7���Q�H8���������"��re��A��i���Ypg��N�;P�فJ��V��Yy�\����m���44��B���%�q���=Q�e��Bδ�h�Ԩ$�����H�?�M����b+��b�e��\ 3��,Ǜi�.�ƹ��lLKzDW���82u]�e⾌�E/C��'� �?��)M�Z*ٰ�y�
0�i�����T)�Hajm�׹�.�_@g7qٱ���_V�3,�v:�^|�^J��Z|�@��/ -���|(���+�<��`�>�e�n�����R�0���`O�!�����Pzt%�;�T��Vm𶘔&�o]�4�������p+�
����	�F�dp�I��w��"�=�5�����dTd�G���_<̏	�JU^�gڳ�q>9���m���l�^`��F�Z�v$�U���6��t�A闡1B4�������;�O���z���b��V��[<�O	yܞ�x���
_j����g
�����Y���s�Lų�‣ �f�����	M����VS�FU8�(0Q�+�@�3��������=l�JT��23�=7��~ª�4�,�V;se��"W����9��A���������_�Ժ����,�/��^т���{j��ֽޤ���L��}��L�ɔ��\OΝ����[za�$���G�,	�kM��Abw���ҖƤ��gC:�|r�d���T�!@W��`���H�}���u�2���8K��r�J�Y�Xр\�C��s���L9��,pze3�9�
�V�Ob�I�齴�*��Ϳ�L�9X�B�i��k�=����r�m�N�R�L���`͉w��U�l�0R7?�pCC7���s�eD#��W~��a��m�
� �u)�C�I�v6���s��� !�/��V2z敵Uf��V����2��}�9h�B��A�W����o�:��G�4'{���' ��R,b9L8Y��Ⱦ�l%�������XA�*DH*�i�ᾒ��R��^F{�jzȄ�`=?�0��.ѥӢ�d`-_y�+��HL��Κc��[xG���%����[���'ңx�N�T����꽴t�4�7��4�I�_�u�!�[!�	����La�y��($q�+�͹G�Ǜ8T2+�c'h��NK��n6qhY�����iͣ�g���ú8uz@�7�9�BRfC�&���&auy�)��Ǵ?J���}��T�ަB��� ���(Y���9JF0
��h�3�_�����o��=	~����1*��o�Az�LO�H/�wq�,̻)PQ���V��ht�|���������c��հxo�{4�����UN�5�ޚV6e�d����~�t�.}D���r"
M1��d�/��t�Z��>���7�k�V� �e	�!�u��jς&[���a�Q��W��L-f��U0���7��G!cx�!ÕH�2��z��/
و�5bS����q�Cv�O�T_�$�ɱȨ��3T�8K'���Q��Q�[c�&P���D�sD���ΰ[7�G����[Ȝ���Fw����}Ԩ.Ŗo��b�����>��IF�ɋ�P��'Pw�f�2����e8+�����P���iu���<�)��+C��l�-��Y2�1�#~�Շ�u2l>��M�JL�vX`чm�$+�N]Di]���8E~�aB�`�F)�=���>�7>�w�sRo	�!�墼�_�?��:p�ǽ���-�����g^M96�$=�)j�m�@����0g�0���i�0��O����'8�VcOyX�VL\�ޟ�rj��q�1�n=r�̧G{���r�\P�$�������	T R�xI
�lܯa>G|6<(q_>m�!�{Q1`���N�%��Vϳ{�����2��g�re��i��O2����G���O�I���ަ�y�"���hQ+�H�g0�y�G:����OJ&H�|���ܯ.�0�b=���^�lL�8%�e�t��2�»��%7�z@~$�/�#��yϦٟw%�7���>8�6P@�4� ����!N���Z����XQz����9~Հhn����6���K!�ӆ($�5qz�0�M~sf��P 5�!Æ�n7ACD�����N�1f�r�a��=�{�1}��V��X#�"����a5�����6��9y.
�k�ƚ�<��/U����A0)ϝ�&�z�S�)�t�P1����-�h0�>5|��;G2� ̳��8���e��H��6�+��_����C�q.oF��~����X�@�0:dIW1���Ikߢc_�������,�(]� 65�j�x�5�bӃUw���o~ǣ*i��#ה�@A���8��$���z���G��`���l�:USNQ;��-[�k�bPm⨩�9i�8���_�
�Uģ�̐ƌ� ���f��"�;��|{��|>����[_s7o��bX?�9s������f�dQڠmhB�G�3Eu��ԁ"����N���Z;�*(�(O)��E�B�/����",�{��G��ܲm���$�
B^�D��o\��T?^{G݋v�E_��U�,�B�U����r�G�ӧ=�/��q��v�q����ՏYWs��u	�`Я�9
��Th�������%����ZKcB)�>����uۀ��R\O��m;<�=68�_����
F�n\�h�Y��1���b���gx�T�#S�e�D!K:����.AEnK�k�D�EKŬ��V0�;����ݖ�TE�X�h�Hò�=0S3'���,�@9XĮ�LqA6]B���\�����؂0V7��p�m�O�^Y嵳qm�3tg���uh0�(ۡf�<4w�v�,��KC	D|*~[�c�.�U���i�9�s�U�A��}P΍'��c�֥@�-�C�>x��)fj7;����x��Ƽ��R��2e��)�~�v�'��'��lȤ���������B��)��Wĺ��P��Ǉ�3h���xã�y59�4"/�ڏ=Jhh���
aYNs������G��2�ǘ�#PV���0�&��>��SP�22���Wh���ߐ��WϘ%��Jp���9ɇ��+��}A謎,�'���Lk�v)�jCV��^�h�Ba3�����8\�Q��>[Q<�.�z?� ��6���L���mKOqU��T�� [0���,*�1����(�F���ߌ�w[@��^�����6�;�444�w��kNj\�R�y�V�-�&4q���%\�>�tJ�_F�H�
������aP̱��_��t�)f�(��:�Sb�p���?v:�<�m�jo�Ȣ��o̒aw�:�$�0I���}���~Ѵ��Q��^~ڀ"Ƀ\sI ��#�-�ۺ$G!Lw�yEƢ%��o6Z����%�G
�f<
�G��: �N'��������V�E<�K�ޱ�|��5L��k$O��r��3������#. ��&��q����]�sY�:�ǜ�{�:9�P��Qi�;�ld�s �xޞŻ�����]�FPâ��b�c!�$� �g��șʹJ�Q�P ��\���DX�+ٌ�c��P���
t�A�X�_�ƌ(��E�!��@��:�hw%�[ɱ�L��O8Cߎs���`�'=��4���?��o�S�Wh��,�7B��g9�y׏�y�{��LÄ�$7�n��34��ep��E����W���H{�o�T=�v�iZ{|�^���H����h��O�cr�H�/6v����cͷ*�ƙ�<�ӓ(��\4�ۍ����-B��>+Z��rz�DȧV�p�'dŧ��,pH��g_�	l�W��Q�%y3Ǻ�@����`�y:�bU�5%�der/���M�@٭�!2K��=�1|bYk�`�-}����(��\աe�yQ���BPv;p��n��P|�-q�f�i5U l��{���ǂbD��&�⽐��mB\��4�p�R���su~F������vMU���g@9^�1���P�(`��(��j�c;���戗�woo�,��[O�{a%�r��%���i�5��"Z[�j6�Z/`�^����=�~=+Z�ۉ��X�9"PS J1g��E ����9N����5����:�z"^h��E�^�r��Iq[cᥨw���yU�He�l�*�ǔ��b�)�G��jX��2�b�&h@(�sN<W)A��b/@y�|qg��j*0�_&VU7�`��ns��_�f�9�?�4��6�u=��Ҝ�@��,]�8|����M��]}t%�|j�'�T�ր1�������z��W��'�s�GvzV�Q0oF�<��^`���A�r0>��.�DL��@��j+�����O��h�t���6<u1^qщ��ldK&������ŝ#p������>^�e�*O��#�Uvwh/���H5�Ҧ���L���d6
���g�YH����o �c�ʫ�ϽbшM9@��mi�(�;q.����h*:v�i���H��N��s�{E2�+���[rI������J��O�ƀI`�(6�"��B{��L�>�~�6OV���YS'L���.|f���$9LwJ��D��f��&���9'��i+:�5t�{qY�(g�C��#���_�B�=�kAE��׉�zf�N�C��_;q"{�#.�D���1��V�[d�g?P�
wL��O'��r��h޳����ػ5b24r�l�W�SL#��~xn�b�v�^�P��bUe <�z�~�㕕��B2�L
��0׉�D��/�L�%��Y�3���H%%���J��U�ov�&?a��!�ȮQ5기@G�>t�ԃd�
s�
�����k��&��V�\�� 2m�}�Ď�LJ���=��QNl��<�Y���0.qY�/Pk�Q�2W@�����C�'u��"�#�e�2��Z7T�)�����^�❈6�F�B�9g*��͸����֑�8�<����uY�B� V�]%�U8>yl�5��/S5�[��DU��wг�X����8��?�8(�Ү�,��t��(!	*�$����.�976�6O!��TB]J���͵` Q^m+2��������j,�5�2�v.NywW2�օ��N����"��>�W��S�0ҷk�`�piA�Z�p&�A'�`�t~��@�Ὄ>dS��ƾ��QR
�x ��/]���"�E����= �<=����{��I,��*��� ��*�ˤ���0�{z%`����>ԋ��E1?)ɿp�S@Qā1mu��Cg��U�J�$[hY���n�S��b�hi���1k��s�_A�Z�w}p7�[�sp�i��i�2�} ��\$����0��-��+�?���<�|Y�r�1o%��d�U�z����Q3���g�.��OC/�U�*i�H�#�!��^���E�2����-'w(U�A	2��Ӭ�}��b)}A�o�����JV��=$DyU�U�����({urm|#W����L��O
[`uVA�<�����TU-�N�ڈoC�eJ�(c��q���+�Gю��e@�G���"��}7sIp�`�&��pb���B�q�y������/�!ȹ�+BY�:L]�d�߳
��2am���.�-p���zf �χ^�.��Ⱦ
w�t�oҬ�ϸ�ݻ�36#"��v�C/��P`��W3�n����gp��Ʈ^)w��HPT����&2��#�0�g�y����2�%�
|�T�.����P�b����Rȝ-Cqc�.�
J�`@$���-5�	��a�56?^��]t�����8
S
RO������&9�_��J^5�4J�]0�A�r�Wi���������k��7�be��(59��C ˉh �[I�x����'K����qsK�x�:t�I����������<>�2�J*�,��,��5%r�� ��xJ��t��;[}���çVWJ���5"
6�p�^#�"j���Q�V� {��]a�A��z��,	ia9��G)�%��ų�с^�V����ٷH*��`V�,AB�O�:�Դ֋�/f�f3��8n�-2���#�#C=��0!5�N��r�w�ī�k�$�|��Ӽ�B��?
�{�y�ca��tX�O�%6�Ah,7�c��:)R'�������9�6��$��*�,��縑�+�b��_M���"k7�@^ޣ
3Iaa�wD�����������%�N�x{�J���Y�6E�(ek�3��[�J���Rٛ �9ڲOI.�j&�Iw "�%�@/& ���B�{ +�ݓ�4ܐt�WS�&��<��pId?;U;m�g���R�3��Q�>�=&�g«.Z^pr\4p��>���*�H �k������e6jS1���W��2u%�e�i��V�U���]�֋�樐������
	@\��F�L�b��4y['�C�+i<�G���vR�Bx�B���蚺��4�p	�)���6O�-�2I;��?���r��FP��X�S$���G��3N�~�'�2jdnL���yU�iJ���.M�dlj-"�,��k[dR�5��0���˲��zy��e-�n�P�=�|吵Wӕ�<T��9�d��q�L���\��ֿ0[������}݋r{���0� �WS�#�22�z�h��x�� !���#M���#!�:a�j�^@XB�%�8�q�)Ի{�13i�:��K��rˤ�iG�����w��N�$o �#p���C���>x�½�<ܫ&��p��I�v�BH��'����~ؿl[Q�x ������+����@׸j%��H�� zs�k	0M�p6HI}�K�<�n���HX�'�<�f"���Ӗ�|��㐩TX��&K&x��V)j����#��E��Y.g�y�I�p{�t�}D$������"�c����o�� XV�r���H��#���(�C���8%0!�����m�uF2�a����=r
8]+$�4�	1�[���	xX8|n<�`3(O�n��_�'���\���/���r�`E&܂S��e����1vM/�׬
�6X)ZW��m��k��s"k�:�5�pVP��$�(��ꉵ���d� 2yسխ\���UiZ��l]tL�~#� ����Ƃ��Ǹ�ʘ�`Y�(��W��c?�u0[Q�V�*�H��a���Z�ڻ� ������J���z��h�@&&_�ddҔVEe(�k9��.��t4!�+sMN.R�\��v������#���s~[X��¨�v�^�.	�pTE4`hH0�	ׂ��J��E�}��Y"��4�������y4��"�0����'Y)����U	T�聡�,(7g�Pow{ACA�MG��}w9g`���xc��|�G_M[���\s��Z��zү �eF�x�oׇrzC,�~�f����
��q�(Wd:�"��%��Qv.�tC��!M�_���$�Hsqv����uj���_Yz��*�z�5�ɨ�e��|�a�%|0�T3=��f�K����b�r[�S��I�;��R�y��3J���q��D�_!�5�����!��O=�C�)������6?x��Ƚ0�;��8H��L`oU�[��;a���e`}6����=��ۆ#Ć`Ȉ�g ?�ʽ~�ЛF�$���;�o���)X�#�N!����n]��~��U���w���F�8�ă���Չ�CK;�����ߠJ6��r��/�^0��H�˳c��E��9��m!���W���UQ�V*񝕏�T���L�Rl|�rv�̇E��p���w�R�maɺ��*�S�m�6
�NO~2�����"@�J���[�zm���	bӖ�J$bʀ��aoN�:�evܝ�e]��(��?����4�@"-#u	��w��
��p�r�m$�T��)h���_.�B#0u3�E2 �����!��ED�N�G1��	�$�o���嚖�.� :x���1k���ư�S�_{@�!���H�_n�7�Lo�-�5����6E-_}-��XD�X���r��=��5 ��`�T$���i�g�Y�Ώq�V��r�i���T��^u�D"6���7��BaFȘ�$�y���=F�,�L��Qt
�dY��TYř&��N���^$6X����%U��,�҂a��a��jɅ�F�eF�-\^`� ��o�/s��=Uq(uz �`���x��'D'�$�)��
���4iN�B<�I���}8n)�B�˭Dj��^�Q"�B�Z�v�w��������HsF=Q�
.!�Ё���<�֪!n��z3����� �(=����e�Az\[��"`b`X<����R��g}l��#�_M����Y�a`��>�6��x�����w�#�1z�Z�\W�͕�娨�}E�w���yCXpΐ���|^O�}�F�tO������d�T�Vǟ��E���|}DΤ�eä���{.&�Ζ�<�8Q�XNr,}���ga�`�rɵM:��A�(R���+֦+1��&r�����
4yinP��O���(U�)cR
폌ew�@� d�I�v��Fc6�$nP\$�T�g<'kʐ|��DY]B��G�t$�4ͦ�݁�ebf�털b⠚��� ���*�c%ěI7�˻����WS�C5G'c&�.k���E������H�U$�*�h:� Mj�Y�k��!������p�p� ��K�o��u�J�Zk�PF�ͯ`����`�dʟd�IA-�Q��D�+�f���7y�W���ڴ�}���80A��)��9�^�QP���{�+�o���?&�,� 41/����DB<v�<��Z���@�g���6^{U��b�V�!K/�u�D�0m��>��*��NV�����~mJ+�Q:�Y��?o�bҩ5ZG?��d�KD�#�̮����ٵM�lh�-(��9�OBFj���*ܪ,Ѻ��׍r)�*��/�����jV�1�7��Ď�n #�s|b�iǫ��0ܥc��:"��g���qc_maj�\�[�@c�X?7�� ۇ��v�/�-�5�36�(����C���AhU�D=�1���>��g_A�NNk3�H�ጨ5�Z�q���Kx�D�����Q�a����̸͠.���oi��D#y֛6�
�O�F��d�{���I�aF�ȀCu�Cu��2?pȳ>�P(��4�FM��p�f	�zm�%���StZ�kH��D����7����S��l�ϡ;���Q<*ԁI V���4ծkJ��cE��̫u���l�/U�����Y0Qhl��u�l�@����Dl<�c3�h.�x�9jo��њ|�y�՜�)��}��{t��e0i��w��2m5K^yE:�:�r`׌Tᓳ�Kճ���)�(�sm�%�����
�睖ʊ�BxU�V��M�F�A�($�A&%�����#�Q����`&���Py�4-��b�b��+%_���Џ.sN!0�7����t��vsV�yޖ9¾-�p]���2�tu�t��N5��D5��@��*�n�JF�i�>�"����p��(4CW�71�%��bZz �N�zNE�r<x�[aU�٩�A��-��T�\�38�S�x��E�\M&~	-o5M�SHg�6˔���3:�;f�R��lnw����0��*&׼ƺ��x�/��A�[ds�̼�6�!�Qn@�\M�_,�*hY����7��qY$�+E�a�8� IA��M�S�O�j���8#�^���#{!�����o�rp%�;eaA�#<`�"��AE:�W^�~h�?\�N�0�#�~7��i�"��Y#����n����9���T�]+���[���cB@RSP�W�MB*2c�\���4���z���[�3�=8qaSc�J��_^"�d�0��a�*)��&����ݫ�o\wd�#RMC�Pp	S�|�Quз�	9 ��l��y�'����(���_��fY�]0Y��E�R����:�~.��DDH^)/���}�)}Y���:�ud��	Ƃ5tB>N!g��kD� �A�7.s���V6j��)��
j��w`�i�I�[�s��\�br�<� ���m���q�����I���l<��̽u��>޷]�!�k�����$�0�l��<�|Ew��I�����f҉�ˁ�e��5���AD��X��������ݑR�&��O�����A�8���l��_�� Avr,
�@����@˅%��w�~iHeu������`!I`��d1�	Zz�xaic(�ALf�%���,�:���w( X���q�ը~hU��[��\X+��	Ĥg�ѕ@6b{�^j�d3�	�.#���}�,=��v�Đ��*�����`�_�����$�-Z�GYagO��Ʒ�z�l��Q f_�<�0;;��:�7!�
(���l��I`!���w��}�9w�G�io��#e��0w���[�i�d{R*�V�,`���t2V��/�Q��H�i�}#AL�q44YU����-�lf�;�$w���/K�a�?D��6²�>�,��D�Ӊ{�j��=5�);�� ��ۨݮ��4E�P5 26#
�>RH�.�[d��d�im�rY��@v:)�z_߄�m��6�ӗ�ۊCft>��h�)J��!^�.�qi;Y���p\��,���}���$[b$؏�����eu�B`���M4�sX["%z16��7�im�2�'�̯��3�;aI�r�`��:����E�^��p�2�9=�w�A���@*k��k���i(���C����7o���@-�\��*_�R���8C�:5��=b�ֻ��>,-��B�7c�J�Q�8�T�0#sD��!g9���@9A�+ҿ��q2m2�h�5�o��vjЬaB
O����4!l�:∧��i��J
L�XBɞ�U��⢔,�:�(�`*�-OX��q	�Ĩ{�O?AJ�p�1>�)����v��?���G�r��h��Q>C�*��
�`5:a��ČC���[�OE�ָQ�7C_�����E�S��D&X���\��Ѱ�!�� �'5��B7����*�ڼB����gTO�UNP,�9��s���M1�!h	Z^�{���u������V-~�JAP�]�PP�4��&p����F�`���:��D'��i�	&�U;�[$��M��b�/]I�RN#�f�Y�NO��y�d�a���4�f�C����t�C�j\FG�j�b@�s��-u���Jҵ�������f*��93Z3�	-B��@���%��D��q��5����ʴ�?�/�*5ze^'W�����W�l��Zb
B��N.Y�5fk<}xT�M�?)J(⢻��� VN
�з�0�V���N7���9�j0=o"��ӗ��SxKw�����l���;r3�>1��b�}��=�)f{��qB�5��#Z*0*�O������'��&��MB�P�؝�|��iYq��a\������HI�Uq#In8�Z��Ot���ү�����mw�Nn #OTR�N���D?w'�u(?�!��{ԅ�#�I[���zhʐ��1���౥���C'.��X�a�?�.B�!��Ă.�^�@�Pb�"�� nc$���:�jb�M�E�b7����ܟ�8FX����� b�]�N�6��m@p&~�_�=� =��YV�a�����Hm6^n){�&%�u(����mT��	�";|'ƾ&��Q�7��M�
b�j��(_Aw?�K���s�V5ga�7�bV�wj:(3wb���=�tɶ�K@�Ga�I����Z!�(�s\rv��m���?D9}"��W,b���0�~U1&�1j����2?l;�9r�XV~f���h��7�A��jEVz^JT����Y�����[Z+�)w{�&ly�РПc�M�˾�����@E����� ��".��Ei��QQĄnm\�W.����!��Bh���~��5�^�f9d��-���U�=.��g��:���)ɓ�'�|e�AQz�"|�]h�b ڣ��B*�[��G���[�w�*%#X�\O�+�y�2p����ջ���}�̲b�F�\��Ȕ�2�� ��ʒN��	��y^'�>0��9a�H����*Gd8N�=+\�� ^ӥe�i9/V$��8O?T��p�s���A�.�(�'�F��~@��-tDll��ӷ(�B�F�N�;�ǫQ���p���-Cpmt美��d��pn(bH��mW�-@�#
�Pz�Ws��]T�R[dX�a,�b�JN�v�jh�Tx1/I�u'���z���έ�����ڃ���@7x*�>�/�#8���+򯄍wĳ�"ɽPߓ�O/+�/�^_�%�g���BG��U�	���wy�
"T�����)r��0�)�z�� �� /u��p�m?9*Fѱ���]Z���_�� ��5j��P�m5������?A%#h�H;�3�M�)e���v������4���d�J�Bp�����i��$��Yn��7��	�T�� �B-vv�G.�����'�N8��D����W��Wl[x�C��#b;�>$�4�9S<�5E���Pv���y�]��NQ#���BQ8<�s��K�[C���I�R�����i��5|�2�V���>_zd��k��1����L$�p�N�}�X�ټJE�*�I���|�o��[�:�1�tfm5���_Nn�B��!������=�v�%�ZmY�mQ�cj�ZW�-�_�`#��I�C�KW���UE�ktG�VC.��l���q�-��j��N=�i�K֡�{�~ۛ4����B�	�w�UwS!��l㓢d��{�fĮM�4�5Ũ8HU��tÆ��m"Q]t��mT���F�:��\^��NQ��$�d��?�!1���>��*�K��"�����d�L�zEpשc(�|fjS����|�����uN�m�r��)_!�*Y��R�x���h��gv�ū��N\-��C�Y|�=��y��oQ��lM�A�ѾUgnQ)�B|e�M����b��H��-��x�1�ݲ��OVdJ�5����2��ҁg)���h�E ��8���|�ԙ�ð���0�s�5�&����;��0D��J0��A8�y�^�'&�{��J�}[�?����(:*r .OҰ@���p��������
�	k���ϊ6�|"u��`�>��;-�����-|�ta���7�I� ͹pL�q�g'�4�u�.&�/��W&j��6$�Mo��zX��8w3eDa\��C�[�e��G�Gn�bNmL�l2l
$�����3J�������z�h^o\�4��y����a%�47tn���c������u�I^.a��NqR��l���j��YZ/���|�d��\u�J�����5�S���$t��
�ة��.�:�m)ء�j�y|�WZVDyN�$��t�,q�<;��+�4s��:��$+yZ�p[�	�:l�yY���-��-<�xq�/�a}��t�lzq��}�W�^�V�Lv��Y���H����e�� ��޺O�w"T䱢�]ZE�\E�4��l5����ѬqEK\,	����w���6 ��MAXO�4���SE�8<�?a'e%J���μ@<�i� �����z�Dz0D�GęY|����%�����������	�pҪ̨�~�.Joh7Z][���%���p9�f��H�Z�ov��`����3y.=ɂ���L��*/�s֜���O�+���@j8-�e��`�$�4PNk6��Ԁ�Ma��MӴUݞ��.uH�CX���P���欳�{����y��7]��GSa�V�Vbf*G�nȩ��^�<Q.D� �+7k��\.P`7=866$Ln�ܤ֡е+1J��M%S��5}y�L��U;J�y9�յ��"u
��gƪ���m���@�U�]{H�����k���ǐ�!�0l�P1�D b��RJ��)q��@���Nv��fӥ!&W�o�!l�V�ɸۗi��2�!�2Q�/�2�.���GH4�x4i7��m��^7ړ�S�A��SI������=
uQ�r���!(qQVfǠ~犉��\���A`2�h�*�W)ӧ�k|���"��-�_�U�ۨU�B��h'�8LQ���ɘ��J��ԘIѧ�>�غ��>x�_{�z�K8��;�(JDXW��H,t�9_vp���"�4���VA�?e	/$Eb��{���\���c2�<o����xނE��@D;$�Ur���6U�6����IC�m�HACƯx	�B�� eǣz��J.�֯���O��;s���F=���YLJ�^c��@�Xd�������c1���uc�����_�6YB�f[ e�_��taew�`/|0���|��H�@h�ԉ⎚=�t�Yj�[������k�\�:���a�%���)��ҋ$�`��,Č�ߩv�����]S�x0�*]�m
 ��rj����D�ڄ�u�J��_ �P��-ya��Zܫ���IӴc��v��o�u��/B;]�����崼�0��4�؉0b�Xq"I�zLN��*jT��j����t��)!O��{�#N�%�_�.�C��7��e. ���t�JȌ��<��T�[���o��⊐`_/�r�)�5#Ǽ��9|���I��J �X�uњ�q�&q���U����ň2k\����+�.��̊5Z`� -�,�梊�ymd?�` �8����w�7p�U�򬆃�c�X{�wfH��wa"kK��3y�	ӑ�p��=��U�5T�1[Ƹy��~D�L����d��J��-A����;}I[E)�AƟ��_wE����!i��3�b�ɠ���x`"�T���}��~��Yz6�H�"��R&����(����S����#�@@$��5��_���K�=���(�jWj��s�����di��D�������8�\��Χ�\�n������e2��ޏL��O��4�`��_$3��8�,�C|�1�ۂ��$�s�v���J����R�'`��ؗ� ��5�W�"N���D�g���ɖ(%�+,��{�����SfY���J��l���n��bf���(~���pԌ�hsoD;0 ��I����1#_@��?�!�/�F�� $���#	�j�=>sPH��*�`�2������9N{J�>P��Y
��A�}�@�˃�s��61�v�Dd���2���ےC0��1��7
�l:��&�QO���6p��� 
�Gك9=A�:@��FP���(�Q㨱G!�H���0AgQ�M�ҖA�u�Z��2���>�Z�:w��G�?4.��눭<��L�,��NE���(%XI'F��ƫ���D�zp*?��	O��bDf3�)�G���tn|*��8X2�~���|�^�OB=�#OG�n<:!�'�9����2�#�'�s�41����6�ݜr�Z�a~�ˆ1�?��b����w#;H���<��a�$�6��ʉ�CEق#����?���`���N��k�^w����,��YR��t|�����S�k�E��cdcϮa6w���Z�I���5S���4��T��������(F�V�yMZ�A���ҙ�P�(������^�m�����5���@�*���D3m���GMWt�$��}������ը4�׾M{�����CR�?u=x��n��7�r�Nh�G!m;�5������{I�"*i�T�o#��wj�>g���6CJ�*]�<�Db'U%<,�!MvNa��^X�k�=+�"��P�YA	�克�"�_F��("��YJ�8CBO�y9�b�@&ܰ��
0��y�������sHaC��֗���#�IeM�1�y}:I���m��BE� i,���蟐Ъ9�@���4T�|3��L��	��+T�*C��X�����&���V�l��q�>tl�gk2�#Up^םB�{�.b�b��v��������\�����{ɾɡ�Zan~�F���[���#@�,?%�e6�1��{װ��N�=���+�o�
�>���禚�%�����Xƚ��ِ.�(��d�����*$K��tj�`J|��"4����p�Ľ�b� N���p	���^,��`�E��2��-�f�ո%:�O��i� ��W�E���6Suo��}��:�õ����x��/Cg��зՅNK���c�$�	5�`�P�}Yql�>��!	��LfΚ�n6����N5^��5�W/���8��ٓ�?0L�rY�0��7;^0�î��u���b��"���?y�%��&"м^i����Y˹6.Lh:w�9FŽ�/�W�PֳD�Ͻ�C��r*�|���P��(k߁=�P"�*i>��@|��+�n��^�<��ȍk*O�]5���ZD�{0O���'Ɛ�4v%�G%*|���.�Ȗ�6Z`,�愨�lD0I�B�Oǿ�p����xmi��r-`@~��(�IۤjiW��,�"�H3D�_V*c�Oo���#TqdAiq�ƹ�j�!�f��r�{<c��(�J'� �ע�]�eY�T�e���������S��[I~�eX�K�D��mT	ݛX{M���}�c} �*���/��,;?�]�ŀue��l5c۽���n�u�3�� bHe�r-���TE�:�����yF�a���kr����N*G6f:��<��Qs��so�Wp=�b�cOE�0�����]{�[S�+S��ak��\*��,FJ3p0#VI�^�0�6qT����4��1�2��B��.�f�6F{B�~jLhp\;H�#�^�Q�`��Ģ�ћuӥ�����Y�b5t9�� &	����2d��6���<����½{R>�䡿�xco�v:���]P�<�!�+����Ѝ���j�h6y�Z��{��Pn�L�*�S�S�ߏ��]߄�_�$n�+K�d��Ѓj�I�صR�z���jVc�l�	�UF��cA=>L��Jl�ۀ �h�����G-�Q����+�WN����#�fq��Q���>�{ҝi�)Q1k�����:/�ҕ1����6�ʩ=#h����s?lN���;k9y��v�_�v��7�*��	j��n����"��6��b�f~�S��-�����Pt�TL#���]m ��;��5y�&n2�ZdIÍ�V�����Ox%�� ?���2@�r�>^ҕ	��α���&��&�U�;��oZ�����٨�n���L���GSɚ�XF�_�]o�k�MYrj���&Ώ ]�Ϋ�VqjJ�I�f��[q�;P�mT\p\�a���C��z%ʇ��C������S� �>c������#������>d���AuP0��3Y�ϐlX�c�!�<&;ܾ���!��j���P��B|=Е�`JHGn��p��w�Qq���X5�-�a�n��*�P�:�y�g�fݱ�����`w�O��{*X���j�̋f��Lݦ-$�G�B���3P;�����V�qUlx�.cr���,#9��	G���6*�Q#�&��~nW�ߓz��,==vX�:ڈ�ye^�P��Mީ��β�k���O�,�����n+dz��ʁ5�S��`@�`��2��恧zO�f�B>�N>U
��-�xv��*ugg��z�X^ěڳ���On�<~�Gn�ʠӈ�T�Ѭ�� 8,�	Q}�����I�xn�~�:�Nb��B�m޼���zq���\p<��0&y�1�>�sW����"n��E�e<�-��6dw��N��R�k҃�H�4��L�I���B��:���P��k{���'����'Hڵ�������Ip�lr��I��'$f֟��_�	�4.�^��������ڊ`�=�k��8k��},NE&�Ҏ�L���ҹ�U���Q�z+���Oiө�#-�D�|ׯ]���=Q�u�le�^��6�������D�ްs�O(b$�`�hY��ΜgPh�;���+�&���i]Bzi/:�F��H�qO!$���vv�o�)�o�R����&���zL��j!��79�BlLͨ� �w�o��]�Np!�{�����373������	O׳�ժ��/ߵ�`^�,\ �0h��/�=��L8��]T�
ǭ�㵒��;��7���*�����I��CȰ���d��[��:m)��S���f�h��xE	�Ps�ER�<ym~N����SP����`�����:Yg���1[�+�s��o;�zX�Y�vx��'ë`ޜ9�M�&!����3�hN�ãU�ظ|�E��ğ�#�;O,I�����(o��6b��;�@�����O��T��4�2�6�m�sk�-� �&���raVTX�H4& 	tP����Γ�j>7}�A�+�Q��ߕ���'CB�`3׉�nw�w�\�6#:#�cr�4F�Ե5�&&��A��]����3�Z��5��~k��T����m����|n�a{4�;G|ſC;Q���^�b�u��\�G���A:���О_sx�t�O��N8o����5�gj���%~d�9���8Ų '�\_�xs|(9t����
��+�P{
*6�.)#�n����8������]�$Ct�7{,|�)�$�3��j=�p��(` F�ѫx�&�h�d����c��::��)��=���^0�Df�x�&�~�u�3*u���� �)��N3o�a�!{�T�����K�lұ�Z���9����Cy��07�I���!�L�SeQ# �_��:j�|��vRJ=�7 ��R-d:��k�
��>a&����6%�ᮣ�(�����W����[�����Z�Z�]��q� �~��� �B����{���.\XҜg�pg�s���C/�S(��*�z��(/�jL�J�~��,~�y�q�u�����f��9}"�=��)��O}E\�)��B�8�'!��mV���
F���%A?�X�*NK���t&�TH،���r�Җy@�f�����^-#[ю�/���˗�����Y2���,�F��%n�,Ú!d�gFps)dWZ���Ri(**���|9�#�=�#�j���c�G���0- H۔,5��O����d �bЪ/��Ԛt��cL�/�!|\�u����1 ��X����&�&��)�wd�d&嶌<0���!4¢W�e;`K�z֒H�ր��Q��/��n�w��+���*�q¥�z�\iaW�T�N�[ˡ����Œ��r%��qS�ө��ȿa�=�p-!^��%�C$1��x+���R�{^��R|�^���4X~'m��	K8�_s�(���Â���+���w2✲��e�c}��<�1�u��/�#8"Fr�!��ӻB;�=A�U<ܙ�g+�_�������bm��붗�rx(c�^b��6���SF>8!T.KS�l�-~��*�,>��!"
���.d0B��l���	٩Ը�P�)�������H3o�%������f���hk��>ӱ�_6�)k�X�%����X*s(�h)���X�Ato,�R���4HO� =7Rh��5ۊ��ê`ĵ�c��U�Qy�t`.{M8cJ�r��4{�T�(�������rF�Y1VXY=�@��mA�x��."����O9v���1���|�Ϯ��4[��ti0=���
�Z������k��C��@��a�6H��~YOq�~�<c����(�T�"�
�������Z��tw\<h�I�"�!ki�h�Ҙ?ga�7���'�5r���2U���m��|��*R��SH4�Q<�a�q���P��ͪ)9$vmg����)@�JZ\qׯ�3���j:���D��l �Dq�[5ä/�X\43,e��A!�Ղ*��El��jc!\�D6��a� �@��8�L���Fv�yn�h�e�}x6zy���k[H)
&�aP���|L�Q	Ƀ�E2���0Մ�bO@'G��w }���N�َy�Z{�"n^������Mز]�4�1�L�Ԃ�S�Z �������~:QX$�39��w֡B�R^��Gέ��l��k��;(7�-jl��oBѻ�Sc�$�|����(�������d�З�0Ri�ٓT�e<eU���n�3�$6z�v��(c���`vzǜԇ5uD4���z5\Dz�)���	G�e���oñ>j�7�j+�����|I���1Hk��4R�~�	�>T8�\�x�\���������u�U���f�v��x���h"x�@,�E;~lO$�j�
]����̩�<�Ń�b���htd(���8��r�2��b4�mK���,���w�]���g~��Ol}���L�l"�g�5&t0���⍹��k��$uw�F���ӧ��WM�Ð�~'ɼ��<�IBs��3 o�B*��d��_��oDd��a�䖶�ٹ�k�8�����Kcs�Bj����3h����o~��<Ӝ�XS���/���f�}�X�q5\���wj4�>�dB08�l(l��pBTR5U��+�u/r�E�t�+=gW����ͽ�D�9A,�v�Y��W�/��\K �!r#�V;�X]�Úm��Î�ڦ2g��_&�X�ȁl"#�yt����fdy����to��=��7q_
Ѓ�|Y�Pվ%�w^�i�$�b%d޲���:���?c�J�������d���7�O�z&���Oa�wr�>Q��A���Q@�}�JC�Ǡ�M�5t���?ZRf�(gL�זi�٭�,���R��e�0�x�����< �?�p���:���4,O
�T�U�G����OBE�߬�۞�Q�n������S�E��V�LW��<f6�)I��D���B���������ֈ����(��\̃z�Ė8���۴���.Q+j�7G`�=���j�W��"��K���0���Gw���ͤH�����t� L���B��y����z���)��� ԡJQ��\sW����)Ȯy�^�e5��a�O�^�m����l0��_�c�4s��؆��t���ڣm��ҰpE���7���Nꖉ�V�!��ˍhR�w�)�/������X"+��h��6�|�n+}�+I��9��m�{�o&y��#!�ȬDo>��i�p��n:�ϟŃ���k~��.��	`qAĩĞ��R���+;v�2����#��F�E�F�H_A� �M&Qm�ND/�[,��kxǛ��w������e��=���7O�tdX��3�k��$���w'��)��q@��^�*K�o��ߪn� ���ph�����Fh/�U���m4-~cuFK�${N ށ�[�m\����S�o��S��y% ��ћ��{3�7�T�<+8�3'j�iY�q�B�#��5;����*��,_��>�|�4ǎ�'�<�H��pK��68��O.m����ߨ��*R��Sm���x�H*@%�9�ljItv?,81�0�6z;�^\����#^�@����\���J�_��LX�W�۲��)����\w������� �A��kp�-��xiB�_�C���Ē;X&Q���u�-��dAk�`gvdW�V<J�p�\ϭ�щ#�qp_�>
�zC�
(��L�p;�j}��3Q�ehYo� �܀�M�d��uCa�^��$ÃA�Ǟ�Q;���S\]}�9{�,x����)io�b��t�ö��D� �E���K������d�;+�����X���N1������"�^����}��z�Ru���}2�
�����<v�6��O�1޼|}�ӿ�j�Jl�&^�G�Q;E���#���P�x��̼v�˃�+b�*��Mtt�A�M@���^��7Q���$b��i�흡��G����엽�>�7�\�-�4z��)��I�wķ�x�B��	�Z�he!��wP49�<9Cnx7Y�(���Ő($(�jN�H�;N"��	>�@\�H4��r�c%����F��H��֋-�$P=�޺G�H֐Ͻe�4Y4�ȶI���g[qx����$�) ���&Q����9Wk�G�F��J�����Z+S�����'�\j�>�]�w��~�QuXgj���8]�A��|��� ޙ�@�l�O0b@L�Y�jbų��ic��k�Tl�� |i�	�{$�\�w�}Qء+��O��O[�InT���J҄(V�&y:�q����j�4b��D���؀� A�f�N��a����6�����;��s~w���Z�y��!���T�n�L��S�=�O<��v�#�0z�<{���d� :��[�'ܚ��WLfZpr�˂���Bh3���J?"$������R�\���M�
����?�����:�7��?[в�<W=E���Qҡ��������v�5{�鶧���Իfbo�~����)|E["l{z�e�.9�^Au�n�*#ϛ��ܡ�LXA;��������6-3Y4��,l�7_�Ъ}GW�)0V�J)V�q�w�ZC@!�h8EQu`���HQ|ƴ����6�T˪�$'��GD�:�Xմq+Z�n	����O�]��ʮ��J�t �ڡ>ɸ0���"/0��]$%T��7��t��
#s���4�k
L����դ�)����umJ��=c�?U�PQmL���W���T�t#L���*8y�Z����n�����`N�+�1�����|Q.!���73	�����Ӈ�������P�kꬕ�u���p-p���X�GOM����V���u�W�Ű�Y����lV���^�l�/$(��(SI��i���_��݃�
�-����:z:�E~�����r�7n�[�E�"�Me��z��x�UyW�':�b�~hQZB��ާ�ܟ#MO){���\b�b��Si>�+~��W�	�@�&W��_�������#1�L�)-�s�<qgeV���9̱Xe��Tj�N,�F7$��d~����74#ߟ.�����~�p��uF�z��6�í�Z0�	��HV�מ>��=�y�B
M�m����@�+�	��i�+� ,Ij��M�wd�����A�0��.BLJ0e�%�ho��ߐ���<��D�Q�)���Vc��YF�ŀ'?�R�Egbc ��\��,��'k��J6G��(b�����w��?Y��Ʊ~g�;[�@ʕ7���G��R����)�8O��}�y�o���p o�"g�����ƵLr������w(SO���ݴ��ub�9k��E�ͭR�)����<Q�u?���*a���ޠ�;��|m��k�hh�4~�ÿ#R@�t��T��oҒ��K�h�k��� �C��]ќ����"ՁV@���E��{�/X�Nڭ��_{Z��d����t7�U����? �r��$r�'n���ȤO��|�nzѮo"(�r��rv�ar��+W I����Dڗ0w��.(c�aDP���T}nE���+�ZC�v����ɒ����'�Ϡ~�e ��1�<oh���I_���*[@�軏�5�{��}0�]_�Q�����  .� �0�0'�bk�`h��nEܪ���9!�O���v|�3����0��=�����W2�vg^H/1ѱ�a}o�Բ�i�W=�LV�!��Z��FLa��~�M�b�W�c���I��M;��[�U��C+��(�W\��=s�)x򄮢4�Q�i��E�u�6�ޤ��b�W$�-�zf��Ht���u!�{3Z��:Z�ۚ�q�����Ԧ]�2{�<ON�9�E��ms�Bņ>���������=�9�>�{�-��+l�3���bw�K�_��xq�7�o^ n*�e��}ك9E�y��-4�*݈�׽��#�LH��j��K��]��hF��vy!Z;HhK��m�~C%kQ���D�:��	�{����q�]ś-̶H�	�n=���;[�����vts/#b'a���u�}��9�{NN�Q��76!
A���	T�����O�����5ߵGu��b?�7	����9����ݵ���1����o4�ɀ��U?�}�oL��Q�1���1���q"<M���9��ۘA�C�˱�7�M{X�7uH�[OB��4e����,σCm"\���[ GM�<4j���آ��A%L1�rlZ0�4�j���D1 k��B�#l�t��}�a�(0=h(2���xIF�Mh�Ƒ��i�D$�T�S�rs{�n{m�'��׌����h߼Q\)�	bZ�f�}���6.9�$����v�Њt�Cz�DkN&z~a�"N(��1�ۭ"98E�����Jj�I_�3�H����O�f�{i�D�"�i:�r���`���V?�tt0.�y��j�$0���Z�G�a��6���rg_$.MĨ������<�T�����{_N�"�B>u2�R]�1�d����s�����f��7�O��g� |q�ٝ�����64��9�E����c�D`�a0�2+�N�=�:�z��.��ci�B��bV�<��8�i��G���1�LZ�|cV��}*�U��e.	�{\�◒����:��B��;�*y�����[oR�BE�3���|4���H���%��M�u��x]G5����75%|���˕%(5j!VSd�)*zUJ�Y\�+3����}", ,Ln�s�,�}�tE�v����m������B�ؼ��tK	��	�(��X�{%�����٫�l�dS�pz���5���G��{='��P�h:��lA^��ap\`S��zjg�\����h ��8�M=�-ī���X8P���?��(Nj`��.у�7[M~w�|64���E.�J&���lB��3{�B�wX_%jt�������6����3'p��R�h��4:�Cz�.�<�,E��bn[��Qd��6�9�v��@��\4vA�ɂ��B��,UK`רC�br7��/	���+ű�r7�������.h�+r�Hk�A{�51�d�X�h"����{�+�sL�C�o����r�r����`4 ��H�N�~������*�:^�,�ss�0n��K�0��b_]�y�< ������w-óc��"���p�T� )E�`�u����鬃�wB������db#�:3D�h���ZZ1B\�4�����=���DTv�,� ���m�(����1�ٙ���.���l����
_���jP
�����e�:���f�l���Ƃ��!���6=fTOvL�':|b\�C��R�˸
Hp�sBYB��jjє��D�T�a��eZ&(wc:gm�x�l�ov��z,�d� 3�OY�}V�ߑ�I�9���\wRR��X���k}��Ά@����<�V6u���)a�Q����ix��±�F��;��#��p��;�-�k�.H.�NF���16q��u�A�������Q8�ٞ�������o�M��r�l���$�~Aݗ6���N/jp��i2�(iZ%"h\�l��ry@�%J�-R]����I�&n�[g� �-��{�2A�P��n���n� 	y.9��W! ����4��ĻM�ǈ�w4���/��#�H�rm �l����K��٪Z���ҕj���f�9��������_BM�&"k��|�P<��́,��� �K�"j'5�p0�n���2w��N7��~5�����k�Z$L�I��~t�.�nA	6�9���x�=���2�d�&* .䰹u����9��6�VV����ҽ��8ɐx��,���
ϤmO��H0�"٬��t�p�+rE��b���h��ic�]�%mH!'��;o�*�1zp9�6��]4��LnD�� ���t�'�����'{�L��Xl'>b�v�Ð*d��,��=��_���o��`L1BP��.���#�\�:��N��@B'Y�^��W��c"����~Fj�6�e%*b�̱�0R}���To����16BJ�����u�:���q�P:?����=�IzG1�q��ǶǙcl�ΟZz���4�2m�H,����NY��yަ�Kv��m�k%�F:O׺2hj;�jǩv�����[��_���J��X щ��C��#/��N��񥴚
���cf��	%y�ۢc�ڶwBLE�TM������n���u�a7�w���I��"v�TAzn�HH�}��X�ߵH����cs�,:���әP����=�AU]�x?�� ��24�>�(I_�0���o�����|]����K�9d���(o@�������7LY��gYu�����M'K�4�`A���6=Nh�iz#��7
a(}&�{Q���O.;/#0�.`���K�r@)Q�G�����AhY���lgut�Bpm�c�Ȗ�%IC���3�j&<�sm��"�a�@R٠�X0n��؇�`�f��Y��a����|�������q�0e���h�k�h^�%�=vP7k���������v�B��h��tC���c ҸCj��vw������"�X�I��V�"���U�u�34v�WzШ�70�5,�'��̏��T�_�a?�U���
Ό7���]�>q4y�:1��o�q7�V
��diC��}�J�JЌU��HW���e|�J����V�������øG���a�DU�H�YZ��r�KMj�_��b{��A��vόmY:5y�)��mww�t�Qx$S��������4$��L-2X�i�A���G:W�`�F��[ܶ���;��DGA\M�*�@J7����ڹ�����P����/������J��ݍ�'�O
��=��Q��;N.��������~I�z��tXi�sT��ӪHޒ.5�H¿�]�S������Z�sT�Y�=�EO��C�׳����ol�C�����(�Rnқ��ʼ����]T�f����0�ћ/F����i�~ŊcdX�mrÃ���J��b��AD"r LܸKM}6���B��q!9�|�6aɯt�#{~n;Jz�k�s��'���q�i"����D���w\��UhϜ��
��n����4�-@�3Z�̉0���w����F��ۊ�P��@���(x�-_�D��g��\b1�����c� E0�)LV���0؇�o�
݋.���(�"�Gژ��?`� t�J����r�u��]g��m��BhM�_F�l�-�:J,��l���K[���m)���çp�W�������ܳ���^�>�jҸ&�<��b��ꏊ�L쀊�E;'�_���ۇK�J|��<�z�i�Z���;@شg��ͫEu�1��r(g�+�-��Za
���méP&

G�R�΢�����qO�H�����
�=p�Ⱎ��g�����"��r���?�Pht����|��(�Jڲq��*c���}K���aS�l��$=�0E����Y�: �h&q3���Z���S����Jj/��@��o?�֕��Ȇ1��y�%
��G �,����}G��T��X�M
D��|��\��8�à�6Y@|��U|��?�i���q_�k��ت����N��d�S����VE�^}�ك��6XO��TΠ��6 ֗G��mh��eć@����(���P�C�A�<߅�#���6]Ȯ�j[�T�J!S�^N�)�`�j��� Z��N(�AErh����<�yӆ̷-�g,R^�8Q�Z�:�d���q�߸��ANuq>��Շ�[�D9l)p5j��H���kC�CSd�Ì�@0)���5-�/ҼE��'�ٹ:3�D\P��2ܜy�����ӶT��8}�z�qSK����F�u �LAl�q]��``�ŉW���<�rA��?g��iiM��"^ٓ�A$2Y%O���ę=�'յF^+`R����ϱf�aY���0�>�~(��?/���}]j�m$��˱9�,����p4�AL<��y��D��b���~ə���q��y��1#S)*"t�ƣIk"<3)h�蘀��K �Q"�����/� $� l/|Q��9�U���oq�� �b�Ƈ�v���aU.z֒�s�U('�r$~�_l8�)���$��%)Q��A����Ա���
�d&����	c$i�p!,�Nk�)r`Q�,�k�TҽOE��'�ˢ&|��ކ{S��������d�.J7�Q����*��A�|�L�浦�ZU�1̾(
�[��I���>�z�3Hkl�o�' ������k�H�S��?�6��V�ד}'��VYk��o9_cv�!��P����/���-�4��3�f�*2ά��u?�O�;�\o>_��T���W��nwQ��(k���))��~�|�dq�~�>s���-��y���=�~wc��4�.ʝ�$M{�fj�&vDc�fvQe��k��:��i!8`��tO�XH�}�i_s���қ+��r�D������{H��P��ہ���Ui��政	������ԩ*B�3Ճ�-�ݢm>��,�y�CX0�9�m{���{e$�P�Z���%5>|	ϋN˭�ԅ�;U��I1-�'��^�!`��d�RK�ܻ�����u˴�`�,>�dP<@rQ^/�@ٵ��q�)2.�YX���,��u扔��pQ3h�q^�
w��f��H��f�0��k}X#����#���[��_������^�Jx'90͕�s2�Z [�}b��l��"�q��F�6'`�us���!;�F����5�׹�o����>��:��|^b�x��ǜr���J0��q�t����!���)`i� �u��l����?��4���Д��R̎7_�, ��Y
�̫����S3Df�9q~O6A�j�.hI1��`�����V�����0ē&�p�RaFF�)���Z���Q��e@�a�TVN�8�M@u��dm�4��L�Į9�A�(|r���Q1�p��'J?h�>@�ߴ6�?�Q���(�4�y�
n(�i��x��"�f�|M�4)f��6��/MWڰ�Ι�y���/��~���X)*;��bΆr���m��'�5�X[�� �Nr�o���љ��l	��"])z�A	�b��SG(��L+vXk�֑I�aw��d����t��F?:��^����V��1�'�S�&�+�����%|��]4�X�r?y�C���K��.�мYUc���l�9�ɳ�&��ƛ�&�}�&̑��
P�T���"���nҍ��k.q��杴
r�u���w;�*��zR�e���:B�z��KN��#�����,��!t��g;V��iǿMz�)a8៍��_�i|�GO�}GZ�z�E%����?4^&�{���o�^ �7�]7D)w�
 �	�T��N��a!�����YAs��<k�#6S�O؂\�t��A�����>r�l)�0Ey�i����;υ���U��0��vx��V�RޱX�v��J�f�q��  ��_PyP��tB�e��ץ�U9�j�+5a f���E��z�,�O���7jS���%���I�_5�GuƖ
����Yq������4"X��-q?����`. �V��W
�7i�u�`�c7���ϻ���Z`�U:�ۑN��|}����xX���W[�����68���k�Md=�7�F��I�?�w�@�v����j���#�m�KM�8[4�;��A[������∆���U[RL޴,��3��^�V}��>���Y���wy�|�5k�3� ��%�$ ��7�7��`��c3p2\g��"�u
x�G6��I���/��G�^����p�OG�i����mȿ���x��SX%�w/�c��������"'x�j�8�ᗽư��m��؏��L���>�����Ɨ�>g���.����p�knDMޛ��7b�1 ����{��k(��>m}T�jZ��Í��;1A�o-
�FV���"�/�z/�_�����6Ա������fz�A��W� Tw�ڝ��W$�	��'��I��V1��@o���DE3]%DHu�6R-4�=e���]]�K��������*�,�]4ѻ�e�^ط2�����2fbP�\w�[��avH�����������C���?V��烾�b^+[7���=5�����˛��e b�|��a_I�����V-��0�}kY�&1�6\״�x��'I-�����;�8W �-�ݨ��K�FQϔ?'ШT@)g\��6a�p�m^��7M�Wgf�:��'@���f�Y�uD�)��:����r%g�{�13�&5�����n雷I�g��	R������C�VR\�jZS�����X�4vdC���Kޢ��Г��U���Ms����><n� UG@s�Om��Byb�z6\�od_\��f6M�E��W/�X����fA��B��Z�����J��c�0��4�����;�_��A����o�j(�;A��w���*'Z�!�)ގ�9=� ��J �>t��<8�a�",��&�-���8�iK����g��U�l��II�Đ�T�i�B#��!G���I�'�{׍�6��y�`���w�i�L����<5�=�/斳�Uo���!|��75&��ZM�e��*y	�(n�߅,o�F��A�+-䚠�ly_��i��MPP���P�/��В���;�^��bf	�F�i�@����@�8�x�Ur\�th�L�E�9
`�
��4b2��)��t�Α��a� ��X̅����q0�؝?�y����lQ��Zy`�7�H�u�rX)�G��S��4�M@����խA����k]6�BM�U��)�)�������^�hÌ5�\�n��#�X�6� ۄ��.�,��������k)b:�i���Fٙ3�?�[ˇ��a1ݎ����Ҭ��L>�_ a>;O�t����a�y7ʐ�o��զ��_�K�O/.�38���Z�n�u(j�������l���r_�@9��r�
�}��I���p4���c.삥Doe�G2A��-�ˈ�9�
�l��3s_��� :<O�ɗ��f��Op���.'�#�	�9!�C�Æf<�:ZyH~�|����b8B::a��}�H@�j��]�t��"�+��O���U��*ĳ��dV��7p�@�ʽ�oo���<~t�f�L#��-���O����H^��Y�+]��޲�y���~���x�NB�5���K��>W�2��"s@�r��'=�<�a��Sk�vl�Y	=�F��f&!����!��ay+Ƌ����F�R����i\9��Z'WPS4��F|(���'�TiH㧗��7�-�
0�{�M�(ܚi.p�}�Sz�@�iϝ^i����P{1n���N���8��W�H��*x���k�� tJ�`�����*�&Yfvl
2�����	Ҁ��"���f�3��&3x���~e͉�hW[v�]�=p,&��>b= �&.��Ӿ���s).
�M�ME����s����ϓ��b����=1��y��HYp��&U��柼:�w���t��rcp*��J�ϩ�*J@�o�լ��)mE���,يL�P�W�,"g����������8��
��#��`v+Yh�*[{��Ø��P�����G�%�<���y�Pn�hg !�����1xfp�TxIz\�wn-No!͔Gz��l��O �i�;�M1x��D�E}���S�L���ή53.��ޚ6�"S�ݕ�UM�e=�qF����v�+7�/���?��6���
U5�M��p�2$j�Ҕ�s��i&����d|���(���:�$S��"�����vKG6���H	\�gդ ������.Zo�D�L�T�8绘�]�vN͖�����!K�
����,���S�@0��	^7��>/�DI?�����!�/t�$<b��N���v���{Yn�"P�]�g^|g�r@�j�R�o���7_����X.f��Jz�cY8쉋*w�t�D5�k������&O���?��J��\�ᇹ���*H&S�˦�b�8h�Es�ԼC-\Fx:)n��褌�q&���CYPg��He�	�U�d�!�������S�2��i�F���\��k>0̲�A���������~��yzu��͞��A���9�&�J���wM(��O5 ���e�F��&�9[��8���Ags��x�v��n����&�<ᗟ�����7Ƭ�R| �3��>�2�� ���Z��]���״�P���|��B��'Φ�}����mJ;����t��J:�F7̂��-ږ�0�����27��i�?��'Q$���*I�㜂��Ka��4Z4�Дa��ZC�[ˉ/��� i�f�,�(:�$}�� l��M�"Nv�����\8DP���,���ջI��ꩦ������1�/YB�h�7z�[H�9@���g7 ���� bt ����۸-��?Bd����RCc��``>'XU:�\���I�Aw �v��Ze�
o��ht��X�P�E�6n]`�Ç�A)���SHo��ԩ���\�!���ғ�L��T�O�o J�]�'�S��Ƌ��@	���@�S��S���qD�-r�^�DY����r����i'0e�<]���[*<�}�b�p�&�/c3y�9�&/��v���������)[��Q�˚Di�҉qW�&��g��⸐�>1`��%����^TZk~�ūQ�t�X�ā�������(��1!
���硠F$����dZY�u��9(���r���H��5Z6#������.1�~������c��#��� ,��R���k��Bd��V��"�$���FL	n0���p1�%�6�RWb���
�H��u�e��*8c�����Q_�~�M�T� �Jb����,dԁ׺j�o����J.�<��
/A�k%�YZ�i3�5Q���j����$�\=�8V�~b����t�r��W�2L�A��
.A�0���,乘��t���վ!�eʤ�`�xm��m�� ]�$Uk�����S1��I�!W?�/t����P��N�1@GVq��zE�ڳN�Ar˝�������\�9�� ��� 
$��E�����Q�B�B�%����m{J@�7��S�O'TH�O/�Y���{����'�ͦ�,f�p�4�+cª*)����S{t,��C�N���Q�j����LX�n�Ns�Y＾��c�G��'A`Q�[2�>Į����>�|�q1Nf�>u	�@�bYk���b���Z�� h��⨸ci�P��tG_;,�γ�)����R�m����U!��Ν*�:a���@���PEPT�,2�y1]��8�u��o�C��/��b��Oy#AN�m�H�LH��z�����H
& ;�/�~�W�ƫ�)�3E�o�!Ƶ�wDpF�"��_�z��Z��I#����2�ÿ<�VS��-8�J&���Ca�0��k����W�C���Z���*��q7����HH����R�(3����	������<��"�q�:j�P��k�{�����|�s���U���9-$��ܢ+��l������v��A�����K�Tj�i8&�T{yu���rN�X�0��zp2qvS���z��]�˫�����\��_�&o±�s�{��-|�$<�����?��fm4I�J�p���۽�}X�A$ ]���bӀ�n��>�d�w��ї��_�4t��l���0��h��h�4(�eܶ�������D�q�'(Q�A}��zL�a����Ͷ��#)9�+��,�{��P�9�_����]?�5~�P9��A��`�.�y��h�8�3S��g=OL�9Ų�P�����#�:��:�{B'���E�6 �N��ѷ
������x�Z-M�]z�����W�Q�,;Q'�V�.�]I5��tTx��F< G�~�.�k~����؞�`T�Z[ec��ax��^EՇ��Ӌ'Նe�NV�	���:���P���m(��zz�lD�N{�ɉF�L�V<U�y�II���T�Qԕ�@Vj��HO�8쿋�����jV���/a�#�Qj��v�5DM^	�
1a���ϓ=�N�H�x�+UA'b>�����J.'����>U亥�+���8�z�"���="/�>i�^�&���W	co��;+�)�e�m��^�HX���U���Bw/o�wn��u{�>����Th��
u�"�u�J��0G�G�(�[�ۭ4~�L6�>D�k��z�?��m��ϒe??��ڻ�aV/5����5�֢􌘙Ë�H&�N�$&>�����R�n��Y����i������;(*��ro��)�ۣ��0��ϰ�g��%s}��3]G��|fP���u�f�b��SһQ�E�/�'����,8�����'���_�p�fǳQG�WBN}���t�H~(9�s�	 :�Q�t����?�a��*���&����e��z��ʧ�1l���R��y'E?�NM օ�ZK���~�.6w�����Ǥ�#��dً~��|��n�,��A׭.mn׌t=�:����
%q�f�X��t��da��NN=�����6��z���|ȯ�T �1֢0�h��L�E�ۅ6~QS�C(5I"ק"j�`����]���\��h�~%��NV
%�Ɓ4-�)�(�%���:v� u�uh�'ᯨI���Wrre}At�"w�ɠ.��I�}�%Nt�qz�M�����4���W�����zv1/Yr�HP����Q%��OeJ��6U�[b�y���t�(������T� ,.f�Wq�
j���-I�G�b�:{@A�j�>��\nXm���We��Ah�I��^�6X��"id2?W��j3�$Pf���Y�?�/<v'����&��ßs�ą�u��!��s�����#�t7�jE���m`��C��;�#x�V	jm��8�l��'!�������ؐ���#x���)�EG��nx�Н��FA8 �0'�P����"Õ�x�r�]m}�O}%c��.|�5Z� �m����aD� �1r�Ծ�c5�9��9(�p��w��ŕ�ƽ�|���WA]}(�?;O����Ը��iD���W��e��,d��hs����d��gKQ]%�-~~1���ü4R�bNhb�$�Y9r��en���ŏ!��ʞu��e�xOx[����Q��p�[=��B�,��8��&2X��m���%�;w�8If���hi���YҨ*
i@��^9{���ؿ���>mZD��3��C�\����+2�U�ߛ!(,f��P__Q��Q�O�!bӧ�.D��}�j�B	M���s�y�[���$���M���Nj���&�?�Ӻ�?<�w�/\?���۵`Z�+ ��r�q�����d������mX�`�h�]6Š:?K����^�-.`��ɾӶ*)@㔼��d���(Bͳ����i1�!/,��A`���91x��'_��u��[��p~��7r4B�=��A<��s%�d���D�?[uܾ�׀5�AS���vbT���K����5����X�JP'D�^��$��~P\���@�_e��y�������u�C^�)���F�[̌��jY����?���*J�� �;�;��ۛ�}L��_���p������]G�~����������0����Ȫw+�V�V�� Ac�$
��)�����Q5��E<!W����ЙY�G�u�_Mg(E�f_E-��Nd��HVG\/J=\Q�Qjux��n��{���8���mYH`����F���7�w���g��柀8
0�׏h|�0ę�0\kt��̩Zg9կ.��C����xRm��_�<|�Z�$+6��1���׷�O��o���P���(.����4kf�Re���mH����ej`4&�=���*-�Λ��(K.[�D�~�~�/�WZ���eE
��@3�U��[΅$�7���t�\�0 x}t��Xj2�X�S+E��a�堽i��oY��#�#��~���G�֔�'x�>���nW�\���~S�󫗕��0�-���zYg<[�ȵ�k�+n�r���t,&�U��S_~)svy�y%@��ĵgtV#�|�>!#�g�Qv�ſG"�a�۷��et���l\���HN�A�Ph��ǧ��C��JF�@x�J	�����L�_h���3t��`���@����[$�`���&j�
L����/p��c����c���}+����r;�Ү�>�:��eb�z�����/kTc�^��|"(� �����.�eZ�����G���<k0@�)0���֭�9|*�js�SԤ��} i��ԸM����b�>�,���p2�X/�����=��X�lP�q�+� 3�=6	�*A��&e�"eq���蓷��D)�z�f��j��F�t=\��Y��C��e���Mlxc71P:�@M��$�~����rN��X`���@['d�Vq#D`m�D;(I�$7�"^�� Ȑ��
�����nO���:gd�����kԽ2l?>����.�cg1?3�4�-$�"��θ�+�V��͝�������q�����Q�K��p	O3 ��tPh�PD���T���9V��dN��<:����Rl��6aj-]i]S�yyZ`Yݵ�?TnBv�3$���PhQwN����Q���U����--���~�b�'H�m�]4���3f$�O#��r�Qx�5F�[����>!�}/�0�(�R�L��.�Z�tsu2KߩĤLW,�W׉�%�G�f���l��5��*���G��J�S	�o�,Kzh�*Cc>M��,��BB*wU���"� ?��䇍~���;]`y�	�����`��I;h2l������"�M|�����b'	17C��j�_��|�g����W3��>q�l8����I����
ɭ5�Y��A�J偀�g@�,�#��U�?�Gt����/�U���A=�Q�4m+.%��#���L�n_*ǂ�w�U���&	p~-Ӣ��BGy��}֐���Y��y�r��ƿ�Y����[-���6~�D��^������*8�s���F��jd�4 �G�k��*We�H�v9z^�^uR���@--����i�ɰR9�PKk��7l�&�2࿜0��X-�Ω�����ŉ��������@Y��}?�uT e�8��Z,���<H�I�:��X �v;�@��sb�!��G�â�\���r�����Wɩ �ɺ\nd�7Zv\Ch	6�z��cs�a=aG�k��/Ҁ|����Ԛ��+4��G�F[L1���f?������2
�K�A{��~�����ZM��ð�g1�����x���1��u���<������>^m]k�A[���u�K��L#����%���Җ�dӢ���/�m�Ui=�O(�^�����noI��xw�a�q�����׿�z.eH�yWu� Ή�=�41�YE���.���=���<�n��'=y%c�9/�3,�B*#r� F�1*	�.��,ͻG�T�m˭�K]K���N�����;�]�J��t��e�V>�g��ʍ����k�	iV���?�[�����oN�@������c�f����*����j�N"�����c����+Eۇ�G�7k��W�8�*<>k08�}�f��%EwHW�&��n;���~��*P�<y��>����w����R}��DNn�XC��dQ;�H�3��'-TBeB�'􏓵)��b��H��Ej�����b�y�i��J�Y��q����BfY�E��L�L�ȟ*����m�`ۏ�
�eu�S�ߪE׽�龂ʛ�Z�z���r�oapN��y��H"���TQ�Y\��	<	v�\��v��l��� �X��>n��=2L����ĿK���� ���,���q;B9F���w������M��Ţ�y�`ڠ�fū���ʚ�����O��sfDk�b2P������ڕ�����v�e��9�5ḱ�(�3Μe�s*|���d����=G���8�?dw���?4ntR3tV<�蒸ڀ�k�A�`��P�ǈvq>��;�Jʸ�h�{����]�����3c �I~���#gD.O�#�Gf�&��@޷Ad��f;���RQ����`��׼q�e4oP���!����g��		^��m��'���QE�3�Umc���mK����{!�WM�Y;�B^���u�w��ɡ|����HI��>�*��VHfP�(o��x��q�G[e��/-�Z.�4���>U��]�у3�g�]����s9�>�P/�/���� w�N�?��_����ycl+_��-j�����DJ��7�޾f����gc���͙�^q<��ٚ4�F+ٵ̗T�O��}� �Gt4�\↞"��"��k#'�vd[���)?�0�e����c�2���ӭGG#J�;��Eu�K�h��=G��Q�띂�P��	l�#�\��N��n�l�4����Kx��1��1:���<ޫk��-Ġ"�}��a`[O��a�;ؼ�G&M�Y�]��sBl39���Y�#_�[�����U��3VU�',���(_���/���8r��QR6�Nh:�������S�JO�dd+�^>�,~��.�k'�LF֦ ��� 	;�۲���E��,z��Pj��4���K!L`�aD������3�{�4��6܋W��=1L	���/So-���G[�+F�w���]``�&*�L��P�.q�m,;�]q��uI��A �e:���I7�F#�ޟ|^#G5�V�ri�0xξ�����?�b��Nn�N�E�oU�ɮ���|@89�U�����A���7e<��j��U%��˲��IT�R-�j�#����Q)��L���4wc���Qa������;1\�p��Ä9y�	&]��l6�sFS�p���71
�)=8EpP��	��"��A���9��t0��FKx͜��="��w��;�/��e-�D����q=�`ý�,����R 1���^����ǖ=գJZ��W�Vi��ϴK\�����J1�B�&?��`��<�D��)��̼fg�2��g�Y��,*wK]a^��1���M�)������Uߍ�����HbK5?���&�c�F��֘���oHL���`y�U�}aRw[#C�[S~�����M����.�p7���`%��wҍ7%Yꍝ���܆�4�����LD
2����������6F���ʃ.ߍq4芴�n�L��Oqs���<գ�sh�����f5�x��^+�� a�8��I�9A�Y��,�eJw�ޕ#c�Ǔp��Z��5��A\�v1"1�	|%K60V���3��&�"se��To��Wuy��3��v�̛ڪ���DM�?P�L��G������o���0~���f&�7y����cVK��$��Z��;��Z�v������c$�g�+�=��:è��"S��>�<���R�幘��p�[���l�ٓ���1�H`���O��&�[}�S�~�AYۮ)�<�o�I�+�l�aN;4�tS*���m�+��fǤ�K���P$�-U�Iu�#l�џ��$_� p �(�.��4"�]A����Nh1�*��2���0�L��i�%:��-�t��2�?�}�!�Ē�F�q��R`��\��Ged6A�����ǅ1%FlQݢ��������Ym?��q�kè���:aH�+D�|��BB��7�v��
�u���0W�9�CMd�g���"������:��ɚ#&��Ł/�M��c���l�j�����}fL���]<����٣6��9Q9�<L27J��_�H<��j�hsѱ�Q��Ue�j��pjȦ9�Z�k�fV��uel\��;���ս��+3e?]�V��F�6��Z��8�'�{�ppeyفVXJD�~NH>���>��#��!"`WE�'A�η���v%f��(h>�-z�`� �H��Us���u�3ĲH��y5	/x�ZP_@!l88F �(�������5���!C��'���>�&b��2��y��q��a��q_�����M���5�<]���"6�-�j���+󀧯a�G�Ǻ���P��_;�9ub�i��p�i���l,T`�&��,F~��;��	�2ɺkT^�Þ*�H���������1Bv�rէp<p;�����:���¦���S���ܖu�(���9h"� X�W~}��,Ѫ�R�İg�\�`v� ��13�5�v�ؔ�F}&�ˡY�SDO�9d��)�RpW���4��*���%8�.#s�,�k��Q�����,���+���oH�+����6��?�Z��9d�䣬U+a���%h��+}N�b��1����t�,���)��MΟec�C����.�ՠlmk8��^qw
�Ղ��R�������^vR�T>�������)x�B�~�n58M���g�۵d����>��	I*�":�dWC3���0���h(�#d'r��lkPC6��:]'qK�F{��鹬Bq��8�֬B�N:�g�x�=0��WU8�o�^HOj���5 ap������h� @k�� ��"���:f�t>�Z��rw��_�k�qy��� ��#~��<J���s�G��7��8ukR�H@X6���m5������gC'�X��Utv��@F��LZ#y��d���Vω�O�]�Q-�����`�#V�Wr�X;�,��T#%of�8Ǣ��;�op�������f�j���>�#7cz�9 �u��;d�J�eBN����o�T��ԧ��YD`��U����~[�<h�4�\w����V>iX�EȻc�$�l:k�A�	%�_w�DӞ�  �+п-�y�>	�Zk����5L8�ί]aj�4��.��^e��_ㆢ_7-ne��D]���|��y,V���.���/���3�ő�V7?+a/��*l�56�Y5F�H���ɉ������Z���e�>���ئ٦S�0m����aĀ�×&H��G ����E��)Ž���O�~��bn��UO�`�����8��������D��6 8�S��ra^ߔ��^xAB��)��.���ޒ)@|Ǖ����hY�w߿�]p�6�bȭ^���s! sVe����:�vz�w�r�D*���&�����G�Eg���
�.���T�}�Kࠎn�u����sr`�
%`�A"�	�Xe��}�p�&�,j�ڥ?�əW�J"��wEbq؏����<�8ϛ �˂��#8�-c�a��ww ?.(F�D/�U����
�y�� �v<�)��r�N ~�W�k��~�*�����-l�k^9ƶ*�-p�޳Ԧ׹u��k~6����h�g-��u3���k��i�o�O������a[�uUI���E8�B��ֳD`: d>��Sc�a�6��u�$�J.��]�/� ��,o�\�7ME!ԑ����7�G$:�]��j*�ϲ�_9��k�U�8���D��ȭe��@ z�? 3�E�����S�R�sk:��.*�}���Q����d�=`-��� Sv{�^�E*f<,i�g�i�6#�fx�[8���L���L؄�-�5,�=��T�Y��#��s��a�.9����:Rח!��p�W�[�9��3��ΕG�)f�a����K����Aɕ��ޛѧ8�^G������aoW��s����N�B׉xu�V�+Y�>[!_�aΤ�����յ�߻��&�P������;���zz˻��#��rӺ�I�Y�T�Z�jV1��X��W9������ѽ
��P�v�zK>ULN��ۗ���ř�uP���{4!�"g���ܡ�q����j��H^#ҝ�v��Q�L� ^@�qa穻\�uiaV:T��!���3�H:Ҝ�*:H[k��yd��]jsM6k<#9
^�+����U���{0"�C��{_�C��	�֍`��F�&8�A<��g�$���5�S��[}"�5�Y��u�v�鵥ng^C�|`#����xzK�\�H�q�l���t>����S��܅*� �pd�7Ȱ~C�|~�El�K}�cHRK�0K�i��h�L��B�� ��$������l���qӺ��fdߖ�n�8=���LJNz����Xb�0;���됑��`�2 �f�ND`p�NwI��������'Z��٨\2��o������|F4�bG{��?w`_ke�ej��4q�9�YN��o�����{ꫫ�	�c���L´�	�b�d�J�|Q�3��B������\��m~�i�,Z�PA�-[��)�������}�(O�¯�%��n���6V(�����ـ�Nُ����ZRE
���EHs;T=����>n��N���`IӄM��4�)�;�x�n!�?��/�wZ���e@	�����\_�u �S_]��w9ˢ�%��V��9�0����=�Vy�k�6��DџLS;�֌�<�Tw����q=?��r#�'k�ώ�FH��J j�SR���@�R#��M�ot�I�.��lAvQчY�V��:j��?���K���t8�C��0𡽼�x;�Y���:)V�3܃`#0��1�F��Es089�Ohr����v��\0�{=��(wVJ�﹀uu�IaE����vU�_��!U�������]eS����,�Z���'�2*�/�?;��i��/W	:Q��t6���]艝�s���U� K|f�
{Pwm� �/��8RY������S�%�Pb��P��|p�i�Cu؞�ߵA����|���D��Y���C'�i(:@���� �_�k�����W�q~Y����gx�FˬWC��㜉?Gί0���zm�/�27�c�_NXB;���	(ex��qt,K?���_�u5�WQ�W��6%�
fR��i���źu_X}�އ�y�^I*�$RALlM���T���o��&le��.L�֋����S3�.K ���0<c2�}���[N�a�9ʸ���Pi�6�~f�zm׏a�����,	'�N����q��*~���1>Y�� T-)����:�'�����-��I-S���<Jf�P��Qc�|i��[�R�j��*�dm�07'�6���\�;걜P=�YfR���R/�	�P�Պ���ė��\�xRQ�w3ʒ�r�L\o�����sw�Ǥ�0Aj�!�W����w<}Vԗ��o�zA^�&x퇗_�@z	��:�oE�|M�q5b$�d
�?,��R3�E��0
��2���u�1A��T7nzgq�+����ƾ����<|{+��,=1���(���c�x0~�r��G�S�ϩ��$��	*��U
tڰݏ&�,8��-rT;&t`C��v>��|b3g�}��K�v�/��q��&��"���;�n3c2�"J�ؚ�a�ر.��V{f��K�p٘E�Y�]G%�'�n�p)��
K�(K("��º%C�-��25"|8�G���c�F,����{�H�o�]�
�V�����M��]� �
\���:�+;���[�WF �btgW���7����z�3�2�˛���#tȩ�R4q�x��K�t���C��ϳ+�����U'�>�(���#���\�C�)��@OK����/����nv�&d�O/0�0��h�G�a��l�x��̾�'=jASxEH�vz�0:����x�0E��!�m��8K�k�t�=o�7��s!f���2�*�D�#J"r,�G�'c5ٞ2O���"��*��g�s;/!�bJ�a��s�]���~[�[�� 2�	�2hnB�׊��G�J�ߊ���"v��w��[	uy@�̴��Ii'��"��e�����6�$+�r=����R��d�ƭ<���cv�%lO,�v�#��(O�O�d�����e������Ju���nl<cj7�������W�1t��u�����!\�G�ZN�d��?�ɬ����x��=��n/�JAY��8و���D�kY��v��2}�=X�v��^b'8�wPN� ���{����d��;�m��3�A �-B�6$�Q{C��!g�X�/��G�/1�Ϸ��B�T���&:���"#��45�]�W�d[2��}-s��O;��!����r��3����;���qR�T�@�^�.=>�4�o$�N��N�!)��]NG����H��R��,Mګ+&u��Ѿ%�鯖���pq����,'C��C'�9�/������J�B�:pf�C�;���L|�wt�%�����/P�u��)�12y��%jg�
_Y����z� ^��*Sƻ�Mh�Z��	+2�	�k$'�x��٠�C�JۖW�����[`�x*�E��4Ԣ���y�e���#� ����G�T����<��X`���x-�/2�
ev�;♀9}т?CU��^��Q��1о�`l�2&,���bs�� c��v�wۛ}���ݱ.ʹ��N�ٍ�┎r��l*�xWٿ�wT��� ����ò�(�S]3X貙�S)�£ B��zA醱�~�d��H�2��p'#�ۖ_�i����^OO�)���~�p>�Ii��
v�T����A�.zq��.� �f�oKu�w�ɨ��A./pvU�aʯ�a СX�,���J����(�L}�xY����_�<����L�q���Y���aS�?�vv$˚��_�U:v�-�gQ���Ά�b�؋nt�*�ҧ@���&�ା�2���J�V��9N�>��#d�i�K
!�y�>Yz�:��������T1�Zj�Q0�x��2�)��6����]@�	-c<h��{B��9µM8z�N���M��h�7���y�+^�Y���qajQ���y\��L�]�����Y�Z����p{-�3)�X[��Ţgu2�D���a?��R��?��w���I��NHʽY�oaf�q��<�r�?�kZ�3�{�C�K�,4��?s��MrmER����w��[��[���V'��&����7�V�R�ěO��\��̐ow��xU(�N����&��ז�F�Ơ���8�@���&�+�FTW��Me�ʯ�R��vʿYﵤ1��2�X��׳i$0jTL��{�t&7�}al�1z���p �@��hn�s��,����C���E�dH�w"6�;{,�Rn��^/e�i���N�g�_9w�(��RcQ�4���vۋUN��#	83�e3l6����ӭ�hI)���R�B�V�3�\MC�q�bIq*x #s�~�O�#m����BD޸s��#�i��W��4�%�f�ܜp���:��2�^���%;7n�,:���5�b��`F��᣶f��J�j����w����Ȗ0 ��� �)��h�B�ĥ�ܥ�6�+�~��=��ł�b[G�Y��F�غK��N�3�'tZ[���ڔ��
�5�L`^�2�ח'Dc^�z��=ls�!N��O�
m���n�Py��x�&�לּ����"��WCo�Jx;���iC�";�yW�C��G�wT��2�An�R ��ԍ�VE�[v�3{҈1��� �T�0Z��\+��_�ӂ��n٣�@{G���]j*�oV��́$�~�6���e�F(�&�a�5�� pk=���פ(:��u0_��7C?v,ȡF��
='6�I*����no��@�� �|Y��c�e�IY��d�i=�����-k��n{�=��ր�CN��f��}��Z`��\uhb�KkSr�g���4��0��Aʶh���޹'�P5qf� 	�p����-Z+�*�g� 4puv����㳙L������ҟ~'sob�b�(g�^�D�ǖh��O}�)Հ�U=:�	�4���z��/Yw1y����j|[�|��(�U~�%7�Q�X�ա��{^ Etǔ��:DQtzz6hF��mh�� G�9kG]�!�GJ^j��\�(���?�)M]L��U���Aw˄3�ͺH�z_�}D�\u�X9]��RzG^��IQ�<�N0]���]�@��T
Z&�?�c��27����S/g_�(����A���m��+���*,zU���V�G~⣰�-(�>�S�,)����&צM(���1:k���xNo�̎��e*�Qيl��x;<ܳ]Yi�G�u���q��O��ԙ�N�h�Ƨ�\��j����Yw����	�Sa�(�$f���	.��g}�s�-/������c�"T�#�S:Î}��ʴ/�J�Oi�^8�6Y�W�qN���"���3�p�}㵰��`�T���,g�/4�.5��ټI�~����C_&��{�x�QH60����a$��_����������$ss$�����m�cA}@D��w���S�=���&du杪!آ�;`)�{��y�O=Y_Q_G
�[�OYS�>���1Ip�41����^Fl�����=�a�㳀��]a��v6�:b��������+�rf	:2J�U)���2�9�fA��2JDY�|��U���w�{�=phtߊ۬��W�T�!wŹD�����p���}���m��l��q��0lxf@X��,^O��B�'�B����=������L}Ko�	k��X�0�Ob@g�`���aW�B��j?F�.���qf��'��Y���aI�m�cj�7K�]�	�(���L�r�u��'[oM[d�'����귲40�w�x�i�����p��~���D�[[�A(��cv�	;�5��:��Vȿ���2��J+�I�����y��A[��_j���K���S0�I�b�3	�Z�^F��bh���j�e��S��*۠��h �*%>H�,��h^��?��kr�	��G���h��m�RdU~�o�ď���)dw*5<�T�Y��X��n�%��GpЩ�Na,mj���dus{kܦ:F8
/a��iRm����r@ku�
��C2I2�擧��R�0ɫ��큔"8a�h�B���тL��<1/�_�V{8,�8��M��B���:����=Z�J�?{yb�k9�L%�u^%�ښ!<�T��n��2�ax/����KRL[��1(���/���R�"()]�|��
�؅>oN,Z�,���$)�H���B���N���Ў�28��4�-���r�4ٞa�Ζ�%�i�C F�Cά��KJ��,uz��v�WN�f�V�0�iqi�]6�#�?��nN�����q�c�d-��P�&���}�75^��h���
f+�c��/<�I,RYK�� �KX[���ms]��m69�Z!�}�J	��~�m?`2��u�UKo��>�T�����rFi��ي�o��Gvϲ$����;n+w��e�5�2�D��KXd���O�*9�L�[���,|�j��DN������$W���X7�Ѕ�5l�2k�R�;+�'r:��=�[�ޥ5���"��FKR�[���w@���)�,�%�mlβ�,sQy�0�R�H(#K-K��յ�r�������F�q\E��`��Ҳ><g�q�N>}��?A4j����SMwh8v�H� Q�h�K�����7����Tt5k{�}�ľ��6�B��Y�n����T�%u�r���?�bۿ�9=��$�� Df�)'4��8:�n�(���Ac )��rG<�q)o0SJ�p׶�O����us�L�'^��՟&1�qj����>��y�R��~�8�����ɧ夨��Jp���u��'o��y��/�6M���C���r�Uު�C@���O�)L�(��zj;_o{@�$�������Z?�]�R���C:ݩ��FG���L����k��h�O�&:�ϳS���z��x��ܱ�����S�B��b�2?���}����i�*�v��� �{�U�_�4X�+λ {M�dw�e�ό�F%���ߍ���q�C�G��Q����kx�f;�쫯ѵ�j)�G�1�J���U���u�D��>���7�	[�G�LD&����'��6�2�NJ��<쥃d�W�e��-��ky�[ҌM<{^}>��E���@�zV�%���W��}���P�@�/���ÌJP��뎈�6?3��5�n>�3�|C�7Z�P�7��D�����1�]�c���������ƭ����^���]�~ev�Ĉ�.��PælL�v��G��Ý���G�M��u(�����#{������Q'�0���qO�-�Tf�X�O.��iV�,F�O�8�Ճ˱2C��2��L��"�ޖ�$F3D�qT��[y2=�;0���G
n�*�s/�}&,*�b/��+1��T!Q{F�]������\)X�� �M��va��4���C��������n���ĚːjCAq���yEoIe�\اT��DS�\�O4�G�ta<���\�\`8���cy%��{���Ԝ�hΖ]zCa �ʛ���A��C��R�	VNګi@��֚^G�6�Z�Ue�(Z��iC"髸��yFhZ��Dj&�E{,5�<�e���� �=PG�_����}M���K ��H�Ϊkzxŷ��b�H1�0�����7N��E�}C�b�LU!w�G�C3��NU�,b.v�� 6�?��\��x�.^��a�*�n���eJ�f�_+�
�a���&�"-M�.����/2�-W����#lNG�Up�ޭ���ox��zL�SW�;�.������#N�����58P8�����[:&��D��΄ěO]�Ϥ��}�-f���Z��>s�/��|(�i������7.?
��7Sj,��o��ӫ��$� � HMxӊ�Q�E�����-��u�U�Gׂ�ʖQn��z)��-�y7�QY��oYq�g� A���j�@?I���a�Ew/�U�Cq����WЦf[�4���Y�Q+D|���{5 G岪i�C�j�����T%��6qm�G� c罣D�;�wR����9hj��)��$�2z�N��
�j����$����Xo��۲�!��\��Y_0�-��Bԗ{�A��?�R���k�'�~���"�Vߧ���^���R0A�����N��B�{���:4��	Y_\�>X���M�D�K�9j&\���#+�jA��f�a�)s�Z�ZrX�77+�aL
X�:�_@�)kܺTbSn_��(��X�Be`�&�+���vM�:�YE�	 � ��o�����Tt�c�e�ael0E���L1;�w���b��s��'��s���L:��4�޳>E��_a��\z��୚pF�(��LX���d��Na*��̇g��$%�������%�+�����I�fG��8�JIi��M"(�+�V�����:�!Ow��6]��i'���r�pgrc�_�įa��xd8Y���1�m�#�3y��J��1���w��ܾ�ǘ��Yn�z����>^�C���%���b���y-X���) ��Ĵ�7zlʨ<̧t4��Q��jWG�\�SdZ^��������FΏ~�);@m��5G��c]��M�\�z\�Zt�&���sh�����6S��1�:�ܷ��)o(�W�*)de�+��o���㜢��P�U���d�b�ZQp`����;!��c�U4�A�0�,;���^�N韩��`���ʼ��Zy�S�xL�a:e�
�7O�u11,B�0����עfR��9oW۹��F*|ka��Z>���`��45{�h&�-�(�k�U�p}-�����t��a)0�P�)XK�Z�{)��4�F�)��(�WȄ5�f_���5dM�C`z !�R8[0�|6�L��p��	wĒ%����=W�-m2+���&����	�É�-p�o�)��`y��������1 ���T8gn��1.m��ZZ���K����C�~�
�$�at��X��i��|�пMW�Pz6Ã&�y4w�]�k��$d�:藍������:7��>�2��'���a��ne�Dc6Z��R;�]fN��݅Zdlĺ��?�NZO��=���0a�ڗE�B��ڹ�*�Mhj�D:��q#t&m���f"����R�y��z��i�[P]So1"�����v��k��-����K��)N�B�y<RW�a[<�
{'(E!(��LlG�U�[�j~��RV�����Ep�X�1=c��%<��^�*�R��6�|�;<���|*x9ǠK-N��� ��E��6X[h'�K�31�Ͷ�AI��˶�X����ý�OX�F��\�JuzH�(��h�T&�<B���#���n�4���ƶ�=��0q����c���K���Z+�N++�c���t�sr�bC8&{Ddނ\�{t��Z{��=z@�������'oSu�GQ���k�aa��j���z���p�r9xx\V	�8��nLR$q7���b�_mZ��wo�����QE�+���َ�f�g�ebN,��1F#�7��iQ��U��e�Oʫہ�+�Ez
J��#��©�H#��?iWA��T�	�y��ɲNV1({�7m��+�:S��D��}U5�|�%�$̅�mnT�s��>�NR��It�u�zC���
�S�D,t"S���Q�Z? ��'�O��V7��{>��5���Ab��&n�3��aC�Ȟ�|��p��t�9v24�S�����bEta���E�Oω0^o.�*E�UԹi�4�Ku�Z�l��QW�Zny��F��>���t�9��J�I��6�+J�O0ZX�������RV���T��9+*�ZЯg��u��b��^���o�$��)�\�?���T_T��E�ɾ��7��,e���"@>p�J�z��	m~���e.1v<\6}����>s��+�#�TH.�H�6�=X�`�Η�in!�a��G�|WAt`�d�����?����H��myOAJ��|OkF�2UR��xfN��v��0�1'6�8<9���t�| iڬ�i���g���rr����W��T����&����:@`��-��_<�|�4��۸m���@��%]Z�E�1Ξ�p��C��E��z 6D^ |���e���+&0N��2�3��Y���z�w�����?XhzQidodB���d"X�$��=%BL<�Iۚ�h2��k�f+�J�Z }�ࠉ{d�|u���I�0N�v����� ��Pঁ}�)O{���"ƴ��
�1|�#���E�>�s3&˷�T\�5oɩG��X��X���|���c&eK�t��]�F�gE�}d�/_}��T���������n}ԅ�(e�����mls]��7�
��eh����_����*��X�j�-��%T����1���V��/�y��чd̞�����K[p'���T��'[,
6+��d��7�s�K
g����+�-b6���<�P��#=1�����x��U̬�}м�ؒX�`aZE��!���S ��2s���|F�q����Ѯ���I�5(�U6��5�9O%�nT���u�~7Н�~4��T� .�g��$��!/��KBsE�s��3�'D��<^S��;�\���_]z��>�&��i�>�nol2䊶������[L�L�w�>�10Y�).��P�rr�7M6���/;�JH>�����Xd)L����;�$Z��>����4�ܦ��c"�r�k��}���}[S����@�Í-	*�6k��{�'C<]�6a��E�|��hGc�z�Y!t��m�d+��9�m�z���٫��\^r/��bM����Dp��Yۦ��破��q'ط��-IĠ[Ħ���Iܳ���7%���⅋�$f�R����Z[��c�q,6�3e���㤣�f�
�W�,�������J�6㪵u�%���ŀζ������?ٱ戟�ŗC��]~J�n��ܝ�;��yd�v����ܗ�ԥ��
)�i�Z��Yh]<VJW,�e�>p�o����9��okc�y2�8��x��kȧ�N_T妆S�NFpS��߾�@�~n��wje�F��c�����t�_F�O,t�Fh�3�}@�%�X�a�O8�Y8
�����,⃰�8$��e,�r H����%M���]��V��y��ޮ�7 %`BX�;�4i�f����"��=���3W0��|b�E�<�IJ��Nx-̦A�^.SO�1l;�͏�5A��7Z9Beu�;�2�[��}񏫶_������eo6�>�CZ�m��� {�r�@[��n#��C,��h'J;ʇ�>M��a���S��%���\B�c�X�IE������`.>��K�R�3� �ZGA���r=3�ǽ̗�1����n������u��f�*mא;������Եg�B'1����c���PS7�?yZ�KQ�n��b�R���d2%M�h��?5���wYkJ��2p�Z�B��N�&�:�QI�q��C��?�>��jx�M�Z�a�.���:����k��N���D_��Y=�9�P���ʓ��1/��b`��^�����@厅��o�ՊAsnb�ۺ�1=	
Eb���b�N��՞�Ï:�&��^5IdT`H6���_U6ቪƇP؍C!���@&T�onS+�vdr�R���<�2'[˳�w�Hh�D4��d4JA�w1x���[ZT�9S�0V!��h��F���eCPk��[ƫI�N�ɺPAj�S�)���{64�$���kp��IA8�2k�3R��4G�i��/$L�;i��l��m���0�������B�.�>sh
�	�P�5�E���6e�=wȒߎ�x�j=���kM{�+,@��o̴�H@���Q�T�a�ff'�a�|!뽇U\��Kl#sV#eW��jǈ�d{hpB���a�k�#�4/GCJ��+z�b��i�#��hv�h �M��v#sê������V��d�ƌ/E����w#��Y��&\z�~m�E��~vM�/_Xr�u��c���Nq�ڶ�̵��Gq2Y`c����KѰ-�[ }-�+���l���L��Q>'�6]�L%����8¾�s�;3�K�r����@����8�q1n�-
�식��ٜrt�8�(G����������h �E��t I���[γ���#�wÒ��+�x��Zy�;�E�k�H�Cђ4}c��&��AL��Ç���2��Ã�$�� u	�£MD�J�H���P��#e��Z��ڢ��6sGwqm�����b�v�P������è[NԪ��,�m��x���g�h�oO��6�9W��x>T.[N�t�=K��Č�ѻV�����ҭ<��5tY�Z�8�\@w�Q7�*�+C���Yi�YIf1��{�A	��L!m��'B�k����%�E�u'�㲇<J^�-k3��!d��=����0����e|;»޶o]�(x�k�$Z��v�Q�sڨ��=Ӧ����7]���"?�W��X����L��4i5W+@��u�  ѣ��6͵���A�?)
�	J�q�b���� G
�;��)���n���3��tGm_��	x�7l�lз5zr~T�\I$��0��b�:5��SlQ��/�rjь��"�.S��ۀ
v�~�`bg�Q+�g�=�fa=W�!'�k=D����1��>b�O�b�ʬO�Ñ��,�S�ri�{)��A׸�R������F��a
�W��P�J*����e"2�<����>/C+ַP��e��Ү`ĉ�Ι��)�$�э����r�w*��?y�x[��3�, ��m|+b��[��_x��aΊ�p�8�z)�c�D��I��$|��Du���(��������ޘ���E��i�jf�
�V��!���/��|�Yw������PS_����ߙ��)��@�lK��o�[b��(\,���|���CE�pcn����~.�UX)�1�Mqs��xԞ3��V
p�d�����Ʋ�@go�k��vfSGc��Igk�i|+�ʵI�^��b/�����~�[?<�����w>���j���ߪ�mNz�O�GM���H����X�.3J'{��=�Q�R;�Lu俸ò��=�7�Zg�2�8�Z��8��M q"����7�޺j���k�'ǇS\�E�o��ak]��Ć��S�������n'O��1ϙ�D�E0t�k���w0�a�Q{�:O!�(DY;}4��\�hBU�v2�*�$�`\^d!�4[ҕ��&8��S}�V�F 	��L2~	��Ϙ	���Id���o��G�}E��͛b�i'V]��9�H^C���7��Gbٔ;=�][��-�*iǠT2����4����k�n���Z�6�e��k���1��&�P���/�G�@��'�o'����F78�w�`a�n������]�:���{-���Xg����0�=�ge�L�}R�	a񝟈����d�K�hxj��%��)�Ɏ���j�L��A�S���O�{U����s��$	R���*8nUa�c0 �A߾`b�)�yL�rG���p)2���m1B�QqP�@�X�}��*W�-��-@�meN��v{�MMK���L4��0#R;��}����V���z�٣��|Tàޫ�n�a&�յ���In����©��gitPB�gJ�ޢ��<�����_�-��[���l۲cV���BAoE��'�rə3������aM�����/���5[b�g�)/���2���?䏐E꣈:��� �}�툖���Y��'�T]Ϊ��zvWIg���F��Մ5��"5��ή;���-VC�7TC�Ϸ�V?������O�w��b���ٞ��~�0������� "�--��N�|�Z��?����4��ɫ[��i����� �L
��,h]"�
�w�����,Ce����Ì������H:��A�k�;N���[��U�=�u<T���賓���J��i v)��0��Uܲow��$���Ì���=͉$|Rc��Z�li܃���'�8a��k����N�E	�������x_8h"���s�vC��{���� i"ɵPBi�����^@�i�v'�t�F��[�.��<��YV�����T(��3���`�"��PǪ�&V,�0s��ֿ��.�c��6��ʆ�����ؒ�̸+� �گ�
5F�q�x��%ƅD��,q{�fs�gXGU@��R�ۘ :��li�������o�$�ð&IH�V��o�+��Vܒ6���(���X�+7Qe���	���(XX���h雴u8��HÁJB��!vd�g��"��ݐF
E��P��lx�zP�X4`'B6�8�Է��� �Q%ZMY֔���S�M���x���D������9��-�A��8�Ih�67o���u@E�w��;|E �Z��XԄ���c
]�����[�H���\�{�U��6L��V��`��i9\�yR���"�-e;�\�a��T�����bP&O���U}��;�U:h��~� tI􈹟8�V���ߐI��g�T@��\Ux��F�0��F��"%�콣_��ʩ�����0�,�؉o���A�v�0�syX%�	rT  ��G�k�����X����4z�N����X��]�Ds*3л�r�ڎ�=o���ЪG�7V����14j�'K�@ķ�/��<P�o��03��M�7�!%��+�3?�5��7)m��%����e��
�V��g��K��ŧ��"����� �r��7O%A��4�?��Jy���!)m��n$�b6��	�P��R���W����'��2p�߂ߍYv��A0��וMf\��мF�}���1�ۇښ�r�6(���%E{I��(�]U�X;e��7�q��ih��5�R�#�~�ՠۑ��G�Æw�sղ\@:�X����˷̯��1�`xwK��0:d�+�
)-�ӁF�\����&f�%̂����#���[����CFXZe���ˎ+YJЪ��9��Vw��m��ɋ��I������ݗ�E\�X���[�_E,6��9�+�LR�Չ	�UnA_;w;+)}�]�š�/�k��?���}Z��c���S�#��Ԥ�1��L~(���C�r�>-��ĭ�Bc�W��)�3m�Ϡ����o�t�	�	=��u�r�r����?T=_�:EP��5��/!Z�\��l RT�Y�*�V�J��2&���?�ٜ�������?;Pi�H	�Z����7ǌP�Ŕ�k���������)6hb ě�A�H@���o��E�r�)�Zf�$L�)C	e;����w"t�ƹE�������P]�U����/k~�B���4��$	�3L��)���o��gS����B�{��3n�IpһA�f�"�a�{*�Zp���a��ن��T�_"7 ��Z�#)��󍽪��Xְ-x@�G(]{d*����VJ�"Y�F/2  �
��'�2ݖ>�@�j�$�.|��NA�&8��
�gj�:plg��$K��4��5id2.�|�{�	�8k��C�и���v�X3�x�����	 ڻ�Yׁ�X��U�a�Y�S���UKZ�r��d̉���'o�7d�|w��� r���>#���9Xï.������h�"Wak�~�6�O���s=����n���vq��^2���K��k_4(�:ŉCev��|�5J(����.��L��,�NĞ�A⼢p����%�F/��E��m0���{��0pM�n��r6�N�$�7u��z�G`�;����W����'��*�m�
JW���B� c*��g���;-̯�-�Ã�o�v��/�� m��+}�E�8���ǘ�@��c�w*�q1 )�$�V�˗���r��1@�i.�c�Q�U����R�hT�79v�<�P����7�0��п���;�H}>��"�i����%~����
�	8iKb �^��p ����H�ٲ�,�Sn3�z ��'�}z��,��:��fט_ꕋ4>	Z��+�V@4��<�&��w�#��j�H E{IA���3�"�� BA|�,��E��a��q�2��`��� �~尰;J�7�����PZ�-'�����	y��/�։�c�VP�Qc�K������>��l��"Ct�z�b�� j? Y�Uf�>�Rf�4� � \��\��I�b��ܜ���m��3��w����j8�O��6�kay���I/L-*	�_�8����|���L��}�1i6����yĄ���2�����ϹLM�KbCZ0q:��"I(�|��U�Jx-���;�/�tQ)H���|,� `)��n|h�]�9ʬJ\J�+�C&5o���x�JPa��H��C3]��e�x���o���b}h``|:�4�\(��I:��~j�a�W�������v�=�,fFK����q��)R��k�_��:��f���.9խ�(��A�#ůݤ����P���v���͓m�ihKKQA�D�}G����8A{�6L6�Y����Իa�L83���ۏ{5)Qy�XB�gR��m��3]��@vr]�AK�������S?�s�FOd<k����ۂ�]�2g]��*uD�(��������8̭����RԢs!f�D,	4v�������P��*�O,��BET�uۗ���s��G�BIL�l�*�$08��_���D�Y����J%�8)e�߿�D�#��oآ��s̽,6D+�J���Տ_�����C�
{��1&��8��N���Fi* 11J_�}s��Q�R��X���_�SG�Eش@w<}����c�s�V��0�T���@�$�M�sd����i���SZ�&Z@Tf���c����,�:���Q�`ǨA�7nM��#��k����������4��Y$Q���1	���g�Q�~���[x���Tw���	�5��ZZ������qm]C�����! ��Ë��g��h�r�hY���(X�_Z���d��4�*e�Z�m���KۥZ������nY7r�����Q$=�	�	��zǔ���OK�i��j�z��!�?dI?�[�-����;ŏB�`�ۣ?�0�A19L�2�� �$�n7Q�@#W��g,X���.��rr��˷ʰ�*�g�	LzqALژ#�W����q�}_ӫ�mYݔ|��� �<���ch��G{]YR������vV�W/r!�6����i�(�?��
�'�:�v����~���3�^�To�����1�DYn�s��܄=민�MTT�+b��"�Oq�����'{B����g'�I~����|9�c-P�C�Mg�р�6	��^�Y���ոb�w�1��B=�6z	z�}�7o�r�[�yz���PN�t	WY��^ L:��e�����G�����c_8���I��[�,���I������v���v����4Q�w�z���߉S{<1=�b'��#~�)�=5�vrK=+�,�q5�&*!�s�
p��g��R��˹V��Q=æk��N�6G�,�G��{�m~�32萑{��]�#����7���sgj%
��o��0	��f������Ph�e���?l��eߙޗ�:��a{3���iC�#	�u/�힦B���}"]�$�L��L0rD��KA=�6�Qk���c�ש 
��m����b��un�ΪN��2wa��Jjh���������;��q�89U~7��ݾM����q�}C[4��kr�k�TH5��
�f��o���K0�E�Tk�C��s40��Hg����.�I�aG�_Jw�� �5��#��YA�mm��{�w�m鄸����nҊ���]�����T{f��i�'�؎x}vHE�?o�����q�-�!�Q����y/���vy����`����*-w���Z���+��kK��`>Ĉ�N`���B��:QC�AK�j�p$�zI�M_�?a6�p��LauqK\Әrn��RI=3!�$:Y��-/�ޣ�굕a���E�)�n�U���qOQK�/#�Q��_�ND:G�������t0�#�������h8�w�����Vʚ5��-Q0��cԥ`2 � Do�`g�w�v�%��6�����gD�"����"X&YL=k	?�YXV6+��i�Y�>ń]e[ب������["��9�5˱*�2C�Y7a�,��®J�K�^����n�@{lȂ����R�b1��� D2�4�����(ͩ��ʩ�J�w_���
�EZ\�ûGt����8�+�X�}�?Q(qO��{�
��_�zd	�:IG��0*��b����/�̲�Ov1��LC;�w��m�d��6��"9��X����VE-{-;�����<	�ta멏�z��敶9-z�11#?�~/��HZ�����1�x��5�}�@ 'H/�~���R���k����F���Y�5&��s��S�*;�S����"���
�c���ո*,��"*J:a���B�8�64�e��hu �廢�!��^c�t�P�}��#dA����Sr����!3Ӳ�p@���MW$+��P�-���W	�����Zظ�;ؒ���L2��տ��Mط�+p�oQB�� E�Qϱ���<j�>�!��@�#"V��ȭn�!|��T��o��	DC�O��W�d�{�,Ҳ�m[����R�:#eJ1��(׫w3�tɋ���@��������5��N'�K����XQ~�!���`$3-!� Ln�ꈁ��a��F�g?�}W�2]��%��KƲ��'7ѻd�-Jک&	 x3�&��^�Y�\i,��jf�/��]��YX4�8����c���#ǋ�K��=�><��衧fD�9M�x���c_ߜ�uB��N�_��u���-�}����G?Q:�H}U�C&�+ڦ�m�p�I�&�Wʵ�S��W����/ӗ�'��S㣓�kT#Ӆk8�F�3c�X��d�ę�ɮW#	��+����O�@_/&>5�&�eh��w.�: �<��-s��1��O�S��Ǳ����O��C�|o�{�󛉉#�9`	�Q��S�aN��Mm	B�ox�W��`�})��+���T�A���w���q����,g���g���y��\l��0���+�e;u��/�_	���c�2���'�Q���@��ȍ��E��9@�+��gQ�j\�
w���+&�_Vqi�݋0�he�/���5l�����?&�%�=Q�j��w�9�E��E	�4[�����<��n�|� ���X{��X\�6 ،�Y
�iȫv�sa�T��"��>�6a�-z<�K�$�/�:�]1ܝ�����G�W���~V�\!��9z�����h_�ѹ%E���_x��'�V�?��i���<#ȉM�8o
k��r�1D\��
�-S�~�H%�x��f��#�w����i���%~`,���y^�%��HD�!������<����D/Oe��>K�����͵a|a⬒X���mQ����	8q���n��1����i w\H��bD$6���E	=�Qj:V�0�t�.z�ڥ�<���R�8��{���W��`�aꍪ���ՙ&�΁�Ơ
%?#�mq�,-�k ���Z��״̨�@;���u�����<\���`)����r�J�[�q<t��J!�Ej�D��l{�TX�\�D��8���E3�ʿ*������3V�~����4gzݲ����_EPa2ec������+���3�b�l�c�g"s.)��l}�K����#E�>ǚ��/	���,���OtJa��������|�Ӽ�B4���̄��Oxnn���t�e)�9�$,�(������k�T�3�b�~��-4ӆc��h���|d�)F��K�+5no�U|&+Erv�1�+�
8�ٴUx�J�z6k��D^F~󻅁;J��u��[y��O`Q�n�]���?�KႯmG-uN�o>T��_`8�K��hƢp����k��Ԯa�ʰ�¥�Z)!�Øx��yܔy&�D ^��:)-A�;�ڰꖻ�cɁ/FC~~�H����@�c�[�)Ɗ�{�⣕�D��!��^�EG��ؖ�)��h�>����$�ܹo�=�4����,�8/P�-��5� t^�M�a�(Z��+�`�����H��+.�� ��TƁ�	��w���6>�l��dgI&��5j�,(�M��W?f+��u��N�
���(Y�tAX�yQ�%��C����	i��=ct���	#����-&Tl:;���9tt�?܏�TB�,���6�iB{���x5�����ʉ��WJK1�{8�9�C�s�@T�v��O��rU�����W��ġ�K.i�kp����w�/�� ��G;�f�j��ЂJ*H����(��鏸zg�<c�v��	(ޢ� ����:qt�7?5q�E��[����r�4W^1�3�ͼ{�+�K��Ù5v`.��oG�Uq�ʜ����t��@
,��W���l=n��V,f�N�V�SH���_�sr�Ag���kLX9�fݢ�\���m�C{�5���S+*8f�f;�N�A�� ��D����<߫�|����^}SR�O���PZ�4�2�Sh��p��^_�-8OB��MtH����/�%��i5�ܸ�(�UU���[��+�1�H}���Aړ���d��r���aM�zdrp��J=��b'����9�Ỵ���~�����쳈T�=Y(���k��b���7n����?7`�EV��\�u�t�����μt�����Rls��0*��<�+ZI��}ܑNs�¹�v��E2���H��CU�*�˂��
���kCU�;}������xw��O ���	@�>�G�� �s�Bk݈�A�D�>z�.sz+�LLq�T@�wl{v ��b��#���VJ3wᓣEq�Z2WRz8]�|�/�agf�|�C���ᛩ2��c�{�Z@}�� ��sl3���}�?* z�I����X�'N$%ņ-�	(|؅OK�R��Al�=lþo�՛�ӟ\���|�0���JÌc1P;T�gg�C(����e��Ҕ��;[���[Ʋ�HeRq�㠧��/o{%<��;�5�%���գ�u۞��K�f�X=N��<%3��ӅL/�ʮS
n6
���lѻ{w�Xe��W�d��X��cB�g� B,��r�ȴx#�	*��4yb���@P҃Ȏ�j��M��9��J.�Mh�i�G~�y�q�vw�?��,���S�8ࣚ�l1�(�*�����O�-5e���Pl��*��Сn,��:������C��}����2l�3|�<�����C�ҦH.�K����ξ�B�1��e��E���u/s��i�,��o�ߌX����_zU��X��xr���2���]�<���[=���D����5E����}Ex%
97���1+dQ5�~���Apx�I%��e�>�t��x��jbIR��N�<Xih~�#}_��)y���z��ro]$cѝ0@��`�7]���)S��r�g�
/�ݵ7����ԋ!�����W�0*���$@�~L�[w:��\������k��ة�S9j�zla���:��]��� ݞ�So<r�S����$Qr���S�/\���%��2ڰα�[Lcw� � o�C���M�Ek�;d<z�;|���8}������L���[[^S�%$ܵ�0?94l�KR� A�hV�Kz���O�qX�X�
�$Z!��9�4�r9��ޫFsR[�f���*��`��ө)�x��,e{����i��=E�<`A��+U�Ӈ�>H~M�c's�j�MVXT�-3��0��q�֮�8��ʰJ���Hah��wWM��%'td��������G˫�D�������"]��q<Q�}*����bD*>}�7Լ�ag��D|���\[k���<���du L>������i��|�V�h��m�"&��&wE<kh[�r��!��;-C��G��S���R�2@�,����G:��-�[��x�VL^������_����z�!�&z_ou�-������6�LƏ��do�W2�������CB�,��AY�~>HP4��+uE��To�4v.|�?��Ku���1� ����|B�!�쁨�5y?T�l�en�.�ǻ���(Ϩ�D�0�T���|��|w_����nh�Rޫ��5�ٓ����~�õ�g���FzF���VѭJe�֞���o��hhgk� &�X!�7>�Ax��?�ě����c@�:ފi�1:�����^�S"	����h�o�߄~�L�����S�:��<�Lj۽&X���+qa�ZHJ�������D��d�NtR��o�U[�*�����3�(�D���{O�'���-&�9O։jK���k=��L;-��Q���B'p�Ci4�u�����VL��`Ó��@$��v2�&�Es��o!�N	Ra���xD�U<ZKm��9?�cD�*�,��%!CSj�
C�^�כ+��0��xK�����~l��a�@���`�q���)��v8���ǡ�7�\�%�qR�n8N_����`��)\ �C����k.�̉bOs'Q�u��=X���AE/����K�7������#�.70��Q���g��'N�O^ ^WlJ�jĩ�Ib�����a���uI�*���(0�N�dH˄���U����d��Hy ���|h۩�jm���P�Э��_#��)�io��k~���iR��D�����#����P-��N��ܨK�ղ���j�n��+e4��o��ܮ�!��/���!]�j$o���M���bcA��Gȼ �m@5		�`s���1��L�j]�4��a�y3_v���e�g��x�Ba��ܵKg��ID6�ĩ�~ż/}M�!��yFw�6�`x�p�K���"T	�}X˩�F�(���cv��v����8v;h�
%x�X�;���%`"v�	��-�!|�j���V'�܅%"30�w]��dI����8�D�q�-w<Ͳ&�2���K���5	Cv�o��\�A�4��v.pdF�5���^e3�^�.��$#`De�j��(_	�@	�n�?��l���h1�bUƜ�Dl>҂[�wFw��❛���2�w��$�t�Ms�e���q��� ~�J򜨊-�!�(�
8��M�ps�,]�e�K:%k���S'.�Y}�'�����k�I��~�;�U�|�#JɑF�0.Q���Q�8fU���Ś@Ta��f�tS�U,E�;��N���X{d_R����b"Nsuf:�ޖI��h����_��*��.�.!�%0I�5P�]����
;_��_�]m@.���E ��1燨V��+�ho,{��ku��7�o'�=���e�N˞��1��z��}>�N��lP�����ڕ��&{q�L�R֛W��ڤ���%�Ӥϲ�^)��A�/��Qn�k:q�z9������`"��~��9�V���~%�`�D�! �Ch�G!�Z�zգce�g%3�E<p���]����&��Fq���i�t�^�_� Ͼ>õB�_�F�"7ȇ�7��5	�ٷ�߉�FZ���me�!d��;	c�,�W������.���*���t����ۘ?)����	�d�gosk��:Q���Fd@��_�QH�@n�q�K>�+�w�5ڴv1�M�Ť>��?��ܲٱ������oed �V�^/m�`���e�'�#���V��aX�&{8����y�Ғ6S�q{w���i����i{xY ����
�J��-����u�׹�p 6V��}4�Ӱ� C��Ç#��k=<4C%ռw輻~[��%"+�694��ý�dJ9ͬ�3߃���(���ڦ-���5��J��5����4q�I�(~�S�ߌM����TQ��	�1�2[7$�_`|h�U�aF@:
W*�p���)9�F}�ߤ���q+.��n�6����81ygoK��1�i���q�O�6�"�HeǮE�a}��nW�Gr��d+�x.̜]$�[�K8����x8	5��VS��mC���ৌc�"�_H��B�~�"(ڙ�QF�%����[���d�R��[K�F(5�Uvn�@ŏ7!���&\�g�̼���縧�F����;�!޾� �x��5�A &��C0��\\�װX���(�W��M븛[���(�P����ǣ�Bp��[˓���g�BIx���1݂o!|D���H�U-zĹZ~�	�"�0C�)���8i�"/�� ���XH9���T_\�&+��=Ynt�'z�1&&z,[$Qz��P�����Wtա����b�ֽ�K�=�j~^�))�h�յ������/��]+!cmb�Z]_�cz�%��]��M�l��� �:�� 'V����&�t�a ����ք�&����ؖ�I�ӛPs�Õ�D�g�6^�.������z������W�g�p���� /�&L?ׁo0yl ����T܌��1��"K�S��h����\���`ML;Z�3R�~IJD�z���e������A����{��p���{�F�o��]¨�97�O���z��0�'�y�:O�V]��S1(�<���X�~O-�IG�H`�����M���C�Q�� b������DT=��84��H�O��9��S�?��}�3�1�]z_A�d.���4�W\<�-ػ��|�<���k�Z����i�h��Xg��)���L�����;�`��{�>�:Ϫ�_��ˣ��)B�N���*��1�i����Xި���.o��qdۅ:u le���O�/-n�E/�W�
_������)�-���hNY)Ⱪ蓭4t`rohj�,5����]�c�{�gtaB��a�����|]�;��9r�������8�1���,ţ��x{�[�et�1�� W�����Xt�q?���%L������}Ă����!���ݼ���c+Ψ��bH�jDj�C�&�Y�^�c�~�i)��'nGj���2���z�����fb�cEiz}�svɓa%pR�a�{Ɲ�C�sS:�SR�Eu�K�L����"���N���)�U� 6�`����8$\CC�ۈbTڲY�=��vA�'�鳏A�/�3'���a�T���B�j�<e�`�v�vt߮PJ�)���40C�UH�]�EH�e��qa�G�g��*�z!$���ݸ	��N�˶5�Ҿ�,ؙu;(��Ѱ�A����2>�A+NB*�KJp�`���#����W��j�G�yM6���1J�m����~��B���BK��d�jk
�X2�",C����L<RO� �S�� $k+�]�(q�\|��`Ӆ��BSb,%�h$��c������A��ȏ�/ٚ��iA�Z�!h��u�ӓg��R����흇�jB6.�)+���R�����bu<RVBآ6�TD��,�;���5ψ����w������\1)H���I.��&.��+�[��	o����RDI�/�����Ep�~\5���T�uG̥����jQ�>�����Ub+.����v�$��Q8>������j����N��<��֒�W��%aICYǿ X2Ey����g�/`�ʥV�Ԝ�o�{�?�fD-��Ú������,@d�?G�a�����/��M2����i�<�8�����K�-�J�X��P�u͌�9�y�NNn��Çj�G�'�%�e7t|0�!�J�*�[��#8K�q�qS�p��2�%&7g�IGjV�ڮHu���l��y�u�U�+�v߉���Ud�t60k�.�eЬ3����:��G�p�.��㓈�+�4]���-
�J˕���jSA�N�W9�0\H\���yX�$���_��[+Y�MH�;)�io���pt������Q��V�M��XB|;]�G��?`}��w����.��Ե����"��-�$/#b|h'g��h��?�+�����?]�2(f�z��:��IG�4�����L��sg���Ѕ��IS���u�����FuKnw?qd��W�y�/-m��f����nf��gA1�#.2�&��`1���muf��"\�:M��B%���z@���,o��y��iY�����i}�S�֤��E;�'0��(�&��C������J��)�'�Ng�b�d]k���ȝ�]���ȿ&%eeX!�6w�_�0��3�v������OM9�mc�R��'a��4_�����xJfr6ג�ϼ��4�f��N���l�j�4��V�qy�w7��چ�x���m� �1��~爗�uˌq���`����b;6dl��Z���~������$߱^+��D�,�B�Ta�؝L��c�q1��m��G֝=�Z�Za�;q8�=$y��=�>t<�I���[���13h㼃���v��E퓣����� e��3�f|K�U�D�a�hP��x�g�[H���'��ja��^pR�ԣ?c�/
9Y	Jugf%��~�������	'��β��5�����^��l��y8ٞ#;�6�8�W;�����/���fS�I�M�"%o�q�Ӓy�%��&�V�`���nm�|�c8���7̀�DO�3���n���f%*EmV���.n���0�n�PvR���Ŋ�%FBQ�?���	9�?�d y���&�3C�;����gk�n�1diO�����3��=���7,�0�G������	�e��3���N�OC�6��u�J����)4�F0���˒�HG�k&�d-�Y�$���5���1�VVYB��?��!R��kl�5��8�r.�V�;#��r���Y�}6�U��k��;�����s�]�;
��}�P�7c���M�W��ߗ�0@K�r)1!x��"�mӝ�)��g�kt=(���,��l�U�Y ��<�`+�>���־}��@x�ل9o������'w��#\4d�f�Ԙ��CǾϓ����s��X	�`EV~���Qz���=��O��Y��<��<X�5���!�=�3�q/+!��|���W��LW���a����9r�B<���(H\|`�ObaE��߳+Y����	�6Z���[0�"�C��J�c~XZ)�0���im����y
���C�fO��`�6�Y3����*���_>�X����!@7�Ƈ�5��:�l��J+sj������66?,e�с�qbsױGh8庬��6;������� ����μP�	wH��yY�ⰙaAr��}��o��hg�
��«7i���р�כ�W��v��[�\�l���O�lUHN�7g(�ʊ�/�|�&�֭K_�*�_�z��;��B!)`��i;x�t$e?#��x��eP��b�F9�fPo���w��`�S�����w)r�BO�|N, Y ��,dNp��=c�j*ZV*��˺vR1F3T��P��	�,1��(��N����BiJ��`|}�T�|��5�uG��8b`�P����"K똻a.A�$�'0������6Zd�\y��Gp��'I=5W$�_�$^�uq���j�J�Ws�VpXaI�B����,��8f����H���t�[�'�rｼ�݂ˌX��jY���7��;`K��C��yo?b��&���T��+�`�(����y�9` f����������?��ttpm J9AT�D�@���Gs5� ��m'���e�`/֦��6�ť�֞�������D��)8=���vg0Ʋ;z7�T;e�1���e])�>��A�Md�,�t���}<TBS�r�:xZ��m$�6��]z���^�8a�1��[69�̋�t�`m�?$h�O6��i��^7t��J���t��N��@9�Y��n2dTLR]-t/Q�M���#`�T!��V�\�E�R��DA�o݆õU [)w�$�r
3SR�GI�Y��OK�����OiӍ%	<�����R�^)��[d ���4׫՚LI��f�}�)q��4����ݼS����Y&�&���w��B�ph)���yk�S#���S���u�p�f�E �Z��W)�SX�o�f��Z�JT�h�i|��!��u��\�P«�li�ݒ��]\�Qw\Z0G�#�(��������"�vzl)?Ӭ�M&�h�D�V�
a<`r����j�M�"8U��i�E��Q ����:k����4�y�o:�]���Y�˺�!��ݒΜ���<���Q�X/�ڼ�*�E*(q��=;k����m��m�]ww��7� ��y⩿<u����gظ�� P���Ci���`�В����'
s�(M�NW�q/������.�+0��I�_���&���Hd8�P��l�0k{j�t����;0�{�;F��L�'P�X����3'��	fs+Su�� !�-.Y���(m�-OC6Ğ�tp��Y+;;�H ~�@wK��ڔL)F��X�APꎚ�H��f�p�p��τPn:gvF�����+�ZWO?h!�M�
���U Js$�L�+eGw�Аv�"@~�,��d��c���"�����u�G8W=?
���?��>��ׂR�Y5Ah�}�x��/��s0 }�9����8Y ���B�P1�.5U�pP�kB�m���Ր���`���m���F�������n�� � 8$����FS-$I�({g�I��U&����lZ�|�"Y�l�I`*e��#�?�4��㲫�y�X���W/dY��}��,�����Of����6 DgUM����b�Z�!�R�h���*蜖{�d#�&ʎ�
�����"�sڲ�5ͱ�l�
��"�?�K�\�5�)���`���.�>n����p�ɺo%`�@¯@��rd��`~  ,ׁI��y����q޺��[���Zd�:2P�c3T���P�M S�dc�`�W4Ǳ����� ��~-�;��'Qw ��;@uC�i�b�pi���4��N�t�6~m�tH	�K8g�}��Q�o;�;9�8q����Z��D� x��6���p!)㕉�3�SaL�����jh��BYz+ϳ���~�#�_��)#ix��c��)#�U�'�9�7E0"������/�~C�����{&�9>F8¾�Qs�2ⲹ�X#�Dٿ�z��5C&S��Tz�y�	���JO � ��'�D/ @�&A�o�0)v,�9�kEzz7� �ֺ< �η$�K�d�HsDw�=F�.��go�)mPւS�t��NXUc�h��^gh^�r��s�];�XI��Y�ٿ@%2���D<��B��B��ct�>��岃�����Z�(��ݧ�sr*Y[�|*"Yۦ�cy�l%������c8�kQ/�"1�E��5��v��3�Q5[i[)+�R��-B�t���΍�u�+ݼ1
R����O�J�����y����i�/�H��U�b?���-��Փ_j�UJR��b��:����� Cћ-%p��-<L�n���M�!�ǺX��	�����y��܅��ġU����^��ױA��V��ԗ�����QE{���IO��4�]c�ķ����M�\A��B�����,j����iT�}�V4�sX�\������O���@ g�lא[�׾����=��!�D�]P9P["Q]��M�at�0Q��Ş�H�U6����D�XQ�HU�L�~�$w����	�O�J0�Ő2%	�7���_�z���M���qsUg)�eE�PZ������0�XTS��'�GSъ�v��Q� �Xl�L�I����V��j Gw�F���|EJ��ROU���l%!���#������-'`W;[3�7=�[��oH�n�i�)J�(ңX��9
���l�BS�eB��^13��B:zǤ���I�����=KDZ�Mw��RB���0E�������)�mj�b���h��Z�A}7���Er��b�@_Ej��Ŕ���&�������BOx�s�ΰD�`nJ�Qgt��:��qom�"��E��D��%�Afd9oy��|$*`2曑�NG�����$-���j�Ţ0oR�y�qŎp>��i�@/,:��Ғ(�-���V�x�6�F0�����99��Z��1�=Wԉ���;�ÀQ��	6E��6~h�͹;�D�Erٷ\T�L��5˅֮��>�����]v�5D�%��쿷1o���ݶ[���R�gJF� 8趿��RR�I$*��	Ҟ�̤��"f�H�0bgƋ�Ɛu>-�s"^���v:u�ى����kI?*�`��oF)�>Z�Y�H�`�@�:����gn����7I��}�]��y�r#u�J�#����j�_2�c��C�-�����J��Ĺ��Vk���դp�L:B� �}Uc�cx��Q�T�ҶA$hc~?�����O1��Ŭ�u��yx�n �C8&�����9���-���&��������_�UI��&���ԋWP�� f����_w;eʿiy��φ@`{9`�ִ5*y�mu���>�<_����=0�Cf�W"�b�ĸ�|��rB��Z�ՏN����<u��J�G3�ME��m5/0�u���e�RO�^�����.5x�oʆY*dT�/����@!�Y����>mXʑU8�Yrf�ʂ%����1[?�4��;;�/.�?�j�u{���!��m�Q���3�5$�M�/	�Q�ϵ벛����4��ә��̇�V˝�'==��MG,����:.,Fg��8%�e�A�3��&U� �2��ܙ�$�`�9WIT7�e�ŗ�Co��x��[Y�!�D,�Td����+!��-��5�K,Y�`�؇���z��C/�I�6�}�z�ċ"l8,1��S�|)�<dh1M�X��cw�8c�p�u�Q �����`�2�f4\�#�T&�u���f䆾�������+VN,K���r}ݵ-�#��#�!�x�-M�d��0)�՜�h#�D�_���*�s�#���������{4c$�`Y>Y��r�K��Y���=l��/�#�e�4�$���үy�Gn��&�x���JQ�@ܲ�*��/4�rK��r֧�)��.*�u#ioz�3&���>VG��J8��b�w]�ԩw?�{F��#,�>l���+��B�>�ۖV(l�T�����I�c�]N���� I����5U�y9�>V��2��7����������f.e<�������9Q�"��9�s��Eq&�����MN&�?}���G�0Ї�6�4��Vb�^3�ph�2n��;���۾#K%'I��g��縆��,�:~�V|�o,|�{�ϱ�C�7iwZ{$h�i� ?�����6��e�6� $b!%��v]���YkB8��u����Q��n�ɡ^m��	�#�M�y:�bl�R}<f��ZK
	�y���f�`�4>n�>��`!>���)4s7��.RV�^�+C�����l�f鈿[������f��%��ʋ ��K<�B>�(9�#b`?�(>�;��Eʣ�߰�e"�
��-g�����^5�)�̄�yV'f3]>&%�JkK�=�	؟CY�|Y�G��B
A�����GE�ĉ��ڎ1���1Õ�[�G?6�}2�K��m�k��nɇZ6�%T�Z��@�:����C�c*^�ߔ;��*~/:���33��W��r�C��ǯ�*8Bʜ�)�TeU~�-�z��3��	���K�9a�{����?Q~�'��c
��	�B�t�V3�t��t�h%�����uz�R�{sK�AS���+��D�C�"��i��ܸ��X�k��fR� �����*l7ǟ���q�~;���u��`��b�}=������0B#��ZV������	���m�O��6{]IY�[�N��z����:���`��T��,hfNh.������3SϢ0�쏂�i�p�DyP=�9(ي�M���)'QZ���J/�����Ʊ���́�9ݔ�Θ�'tk`�'[��0X0B�k�h�]3���o�Ik'�{�̬�]��J���j�B�ѕ������o����m;mۆ�j�ѐ�ͼ͖tY����#�&�̝N"Z��3,�;���?��۬��P��V��$iU=�D��k��k�L��:O��w<@�4��������s��bE��?+��q@`����l@������qVI�v,I����Є0u�V�0��-�I. chb]3
��Ux���A���EC����~N�s���e�Zt�|&�&��ȃzJ��
|�kuf ��y"js�|���5����YP�<	P�t��"�R�P��YW:utQ��w��~�8�;���}��L6;U�Ağ�Zƨ-�;!um�cǋ�� j:K�e/�w�:&k*�.��?��@�:�1~������``ô�/���Ye���$w�ף��u)�^�M�$G!D�i�1;L'q�MM��jIH����*2���up��g��?���;d�;N�d�YY����2�:������.�
z��da�����g�fRM�x͎����Hʓb�=���Z��gM.�BiD&�8ψC��F����P���Oe������k�.[�I(���aEh�]c�5?3�>��J�I^��wgw����H�<-gQ�cT�?�5")U2 N�����~wE���A�|gY�@��ͱBAV!���.v�t�� 3�� &��C�X.6J|���6):��H��p��s�fe*�3������+���g8�wr4!�R:��C�b�#��K�F��f&Y�J��ed�u�]�ˌk<���ڤx�	�iG��PE�< �y�6o�s$�-s�|Y�C{:H�C���e�X6N����{o2c�7��^���1D],ջ�12�MR[n¥���;���	��7���WwAap��S�r#5���-Da�p����\8�
��5����#߿�XbF�20�v�����ho	mr�������Յf����D9��w����l:��9���M^�i����nS+�%S�+�d*���sPp% 1�j{��ܶ��n��%w�M��,y&������*D���f���Eϔg�z���Gޛ��*�8p)��txdf�nD�f	�G%o/2^c���^���4�͞w��Yy[���J�(�I�c�?rN�m�x��m�����t��<8t�O�f6����K^4������`����K��aP���V�%BYز9O�mG��;b��R�w߬�)��t��6)�����kS��#�Ԛ�c� LA�{e��Z�2�.~���:i<�J��d��v���t��q���5�ht�;X'J�
x�M��p'��x� Zmv�)]��U���X�k,�%!$��;o�`��!aZ��\]W�c��#�@��C@%~�4�
�C�#�F,Q����蘐]��<�Ĕ��BD��!�e;Z�����uR�l������GR�p4��@�,��������)�ͣ�p:�K�Ӆ�^�S�e�B2�F�� TXĳ�Ա`��o��xn}J�
}�)ܛ ���Z�\���\^YU1�Eg�Y{��"t��H&�1���1]].F*b�V'p����ևQJ?o��5b�V��X!NVrА�%D���0�%z���)�9���;u�t���&�3-Rŵ֍������� ������ u��|̿�l�g��Qz�=����l,t�nK?�C���a����p̄?{W�|(�{+yոd0��p����-�?�bl��)=U>���(m�:�q�D����6�{Dp
�B��E����o���4������s��:ڱHv�=��*YY�+Zi?]�ebC�>��V�θ4��m�d��,ݍ�a�.�WO����:�o�Q�Ћ��-������Nv�,[�P��qm��j���>unbMF�Z��A�C����ȶR5��8[����%���B�"r
-[
�Z�s`�h��aw�H������#��H��8���b��́B3��a|�f�v�7��pt2��HC�����Q�2����w��u�Z�B�L4���o��W2������I-�m�҈p�����/�'S[�YT���/�M����I�b:(��;��R��BV^�F�j�;��u��V�toiN@�+\���790s"8�#wHrK�I[��G&�}��r�*���l��,��4n����y�8���\D���Y�gxl�K!ŉ��+�T�k�-�D��ܣ��i����e�)=>4��ܳ|�=O�UX�ʎ�!G��{��I	[��yQ���[�J��+�҆�b
O_g����#�J�/1{�7a�I>��xaZ���y.���s��&b!{�K����̓*�up��0a���Nя���"��E��S��\e��Q����ulX.I��(��b��]�M��G:��j�����Đ����'�SZ�T�u0� _�eCYw���;x�Y|�����!����ʄ{����X!��@M٦��e�
��r�����*��7c���SJ�ʗ�"��t��(����f:����%D���p�G�ÝI�
����xbʰ����M�]E���l������m�X�l�>�q ���\N�X�{.��Q)P�TW��x�h�V"�������6�S��I^�ë-���^ʓا�p�����$�@�����j�(<�c�\Ξ�m&�^C�5����'˗h[*��Qr�vV��A������w���Ց�� ��G'���Ѫ�R�H�G�
~p�^��=%���r�@���:M;Ձ�e��6�t��1�h)�"o�#f�T��w�r��<3�|b�����1�8��+f�̩bǸ_"�������=��G�y:ú�C��d�τ��� ��Q.�h���#��a��S�&�(
��èrl!EE�G~\���]}<論����?3n��+9WM�ZKﯽU8�XU51�:W�@o����C��Y����sL��'���v !��q@X��汔3Ԧ>�ܥ�rY�����$^S�>����α��d�G[W8�.�H@�H��T�+�����PGbS��u�k������5+m4M���\�l/�t3�	q_�"R��|rT��PY�6��k�t��YƤ�����,%�)��J�̆#�y�k���$
3o�ڤ��0�Y�z94���ϊ��t�H��ct#p#��2	Qm�ծ���*(F'�����|��bRE�'�9�.l��x�>��:Y|(RV�g�֩5(�j��V�Jv�TDk�>��,7�{ߑat�^GȔ��"   ��q��%��S��V,� �^fl�ZN����n^�[��W��VlD]6���ׇ���S������u�l%���E���B����t��Ff�EK�ȿ�S$lI�?H?����M�>��ud����^�v@f�.s�f#)�P��z�b�[O] ���{���wD���^�,Ǝ]w=�s�xy\�E=ը��6m�Qh�~�DQ86��P�Xe��B�A�;�|I&o�����Ƣ������W�������)[\���4�C�7W�s��;&Tlz�o��aa��|6~�ͩJ�s�6�>��T��L*PWP��ƶ�UC$�yw���E�C�T�����8$��4��=x\�%���ؔ
X�6/| ��0�(i}U���-�y�U�۷^�MR�*r��E8�g���0���7��H8"L[�w+6z~`8��{|�+E�BP3��Ψl"����wf�Ī�:,YSw���r�����+������j�|`���,�6�58������&�b�ٶ�~�i��p�4D5å��4o��sw��� y���_�J��f̾)'r���+�;��=ޞ[/a�Y?9�m�z`�Ä8�+�xr����N\!�g�D���,K�HL�b�c���Ѭ'�{����,�Y%��	�.���K$��0��^AdQ�T �c_1�P)j�G7��e=ݥQ^��W��n���(p��tg�k�*��\*���z��x�WH%!�+a��X5J���z�ÿ>K�Hl�_gmƅ��9G�=���S�
C������#M\�/w����� ���fC�r���*�05)�V�D����I�ᓬ�@Z"�A"��q��-�%C�F9M����W�:vK��M�MHMzF'�^Ł�I��v��Lg1
�8H�ܻd�45������e��Z�.��c����>o��Z��^�P{�?��B�;T��]	�0��_�7>J}����Ʀ�.�!
"�{=����\^����1�G�:���^�(��C" �D����?^��꽨������ X��X��������N�'P-��<��*G��5A�H��ʚ���}�����L%�F��`��q���e��M	�Ѧ*�����a�g���.JB�ÓKu��Ŏ�Җ�ˤؓ齻/����-JW��k���]��\i��%��J�0�{���`YS��X(/=%E���U�,C�G��M�(jm3����H4�BM�f��6�%���v�l���Ά������C��/�Q8!��Z�ϰ��tg�s��3s�m7�S#ND�nu*�� ��={J���L��kzAsr3qܩ]�S�[�[�fʓ[���P��yY��D|��-f�辤Ӿ4�ur=&��|[�6���2����W��C=���]�l��\��Jv�sĖ�L% ?���g�ا�3i	Y���&�-�)���r����I�,r�C��|����!�AgZ��z��:��S0����D&��yW���;�$�Ω���.,!;�;rTai8�cK[��`V�l��i�Ę �j񩶇��5��7�����UDHt��^r�3������#S�P��'t��6�����Ɛ�1�.�78ޑY�%3W$J�g�Q6|<?�!F���������-H��(pe"߿سe�Q!Ň��T����/���`�ۧ\��@6ZQ��0�h�X�! pn���s$�;��`��7��C��&i�
7�&�>�:m�t���6��&֋JbR��y�����%\׌�\Θ��Ծb��Ч�������6���������aSRzz��|d��TTK���¾A=2��l'���}4����p��5�d���$�[^:�ei��g�^:� �֩�JJe��`�'��P�.R�]i�j�zk�eV���kF�U-����&^���]D>͐=VIa9�&������t,���>�-B��կP��0`eL�>n$��Z���X�� �|Iu8�o�#��82�(nF��G��(���իO��;����eD�b��n�h� V2=�L�2�1O\v=�v�]�#���pc���vm.�1&�/�2Px��w sҮ蝼�����?�W�}��(�9t�bA�w�L���v�������D��>q�c�,�S�w�|rxU��&�Fy�b����@��#j����]^q��|�N�^)�	>��L�D��,��3Tmm�3�s��>Y�����6$-����4�����}M�"��X���A��O���U���B�q�K>Z2|U9$��Ϳ1������v��qRپ� �Qo)�yܱ�ap瞓y��銞�	�(x����s�&�h�z}�
�V̫�
�dW�[[��~�� ��K��7�ҿ�k�'�܄���\�����3�e�T��ŚT�8=�t�G�]y_�^�Ԉ,�O�s͛�S����Պ�ِ���S����^@����.��*��1�*�Y���K�O�D,CU� ������X\�=kE�c����������^\4���z�ח�/5�@�j���vuG�G��$f���|��&�Y�_hS4֙�ܧ��w�׏p��@��YFWMY��.D��J��|g����Pף�y@��nV39�5������_i�T/e�˻�\��m�b�P���bM�Φ�'_���a�*�������W6fӁG"�T���rR�8|��Ѷ{*�^eޜ�ڨ"��E{³�8�����ⲇn|rZI(v7lJ����,YW-����}�ٛ"��ː�<r5�Ξ�|!�ҍ�7g`�*�/7�����Sp�gB�S-���/۾�z��櫔2?
�%���Ԕڰ�9x$�'/��TX����V�X74B7�U�/^k���ٔ㇆���fج���`]be_��f�;�W9u
C�ʿ�Z끙/�A�l��ִ����'�ER�Ɩ����T��ԓO(n����ۯ	��j�}�ƫ	p��92�i1ZI�=�#H�g���r\u( ��K�"qʜ�]�| �+z(�+�uN|�#Qd55� ?s�g�rZ�$�r�6�����	�5G�J�_�d��I��^��r-1�:�~vc�WXXnJ	��k5�K`�@��`̅�,��0���
/�տ�KP�I ��3v��`�`�ޠ>mi�,��\[Q.5 g�)Ou��b����e0�~�R�ؿ��9�s�y~,@Yӥ�3կ�(�Y���z��}�:�Y�lęr�p���!�|N�J�TH�D>�(�~u�Lv(�괫���9̒��߫�P�G=o�7D�	�g�H͔����̽6bN�R��B��B@�n{7�,!�q�57 ;��l�qS�IeFgc+ݛw�� ��HmS`|�,5~.a�?@(S�F���W�/��BU��T��FuB�[��c��3����J\�~Z[.m�lW��d���ZŔ!���Wh}>v��ܮ9\���!��	�x��>��|�������+# ��Hݮ��yݴ���6!z�9ɼ�6��l�F���(��\%#�#��ָ|��R�մA!���&B|�n|o�8��N�y���N�����T�t�}���[/Nau_-��P�Ά�ؽ���̌�iBM[a��L^G�e���N��tK�x�Dģ��Sz��z�g=�U�@���
w����a��'�����fB���.���@}cV�h�@~
%�kk��C �k9�� ���A��󿥤��flI-g���RZX�Q?�[+�S1u���(�@����W%j�^�:A�� >[h\n�&��,Wr���q\av����2<����6t����/]
��2!GK��Je�����3��*�`鶑 ��G�Mp(���yh���{jI�k�:���M�,�����ʏӏ��h��L��,�u�]�ы���t�F�P��=�/���$AJU8�Iz�<�o�� sK�(�Z�0�
���ּl�=vh�	�t��>��b�����Z�7Х-�ax��t%|�_���"0�M���I�ʹ���b��3�%��E�؇��XnE_��[�&OvqB$dI�ş���T��mꐍ} ѩ⦺��B��+
a��x�H�����ꂟ- �}P�7�1�	ln<��Y@�jk+e�G�nW�1ܘ}~)W*^W5��~7��UxH��nŌ�������7�k��Ƶ�����H����&=G!\��Q�Lf,��X5D�!���C�� n\��|�N���^�l�'��4�uI�t�03E_�������dA�#zP�?��&?u��2�&�fvZ��½nωs@lUف[�I���y����qL�M<}.w�=��e�*~߂f�(��̉�5�f� �K���mii�pG��Ǳr�x���˪�K�:�� lh��F������B����%�R
�Ñ�����84|�O���)D[���Iʜzy$]r-F�44B��-��w��r�n�Bk)��@�k�`�� Վ8P���L�ƻ�dy����������6U^wD<�^��Ӟкw���^�1�7S��+��:���)���Ri2bnjأ��1�Љ�:�V�����V�Io�e-��Oa-ע���������[T��Uݦ�ۡ�������
�:'�Rt��t6�SY��z�Iv��,�F���E�W���g7*�Jz���#SϪ��D%��2�k��j�d@��/����	��٠�?c��
.�3��(?JsW���~���[���r'��?�L����Q����έ�AM�k�$�9	ߺ#9�|J��u74%���2�!��4V?��Č���e]�t��� ��z �hiA���&���?�<�e{���2n�|*^y�p���l�7 [ @˞+~���C��4:��w�ߐ�	b�B˶�m�Ǧ؊�\��E�S�wy^��y5��mW���ʎ�����7ˌe�����X}߽
�>uƑ�N�0l��A����KԲ�D<Q�[�{F����߽Yʰ��U0JU�}��F��zM�Sn,q����ӭ�EN7>��z!!Ӆ̗ v#ʥ��~��+�6��KY��D=#A����� ������n<,a
Fb�=��^���]kO3:hD�9���_-=E���i��F�x/Ɓ@2��*c����M������d�Q����7����"R��#������e���S���Ó�x�}�������G�W��&M�26��
q��ks=��;C��!Ƣ��Sb�Pv	J�R	��(-]ȱa��y�L
�w&~;���Ռ�}.��j��dɿ�ZY�*�cyc|PN�f: �r���S�l��+v?����]x|=�/�v�B<��ehZ]�2�	�J�}�t�^��x��	���aA���'sͶM��g3�Q�Ցx�P��9�ۦ�͒��>�U�n��Q&.���^�pȻ��?=ЯRV��N��e5�~�wx6��Q��N���w��¨5iy;Ť��	�!a�X�)s��? -��0�mV�WA>�ʋ�/X��/��]�Nh�K_�Ѷ�H���c��h�Wj�W9��*�-����AY�B%�4��P�Z�����~���?��z�=�_& �f�"fTM?=O�3��W_�u���l_�s��)d�6�f��*P/.�+9�h�jN3�Y���W�WK��<�nL��(B,k
�޼&�Q��KQ�7�sv/�C����:%�+��<�����ʪ;�q���f�ݩ^o3�L0��_Đ,���BV�J��	mu���v#*���c�����.��vkL�G�z��1,	�'*�VMyp�#/E��EbN����P�>�EFFC��k�x��;0
)5)cI���_��:�SB\s�2u7)J"
�k�*�K$�p�4$dnK˶��L:��X�}��
t=�	���r��z\��FEu��G�૛�e��pk ����aUN��d9��:�A����?����_@!��ט�Z���X��yQ�~�J��/���\?���;iu�~�S�)�$����k|��ֺ����|_�XJ�.�q�t�����wa��`�@֚�wkJ�a�;x$�5/1o��:��8��_p�b`���ǈ1���K�u:�`�-d�ƽ�V?WNX2f���-vub��1�M��;�_�%�u��+�l��P&��j�����a���v!�{KUo�WN��µ�2X+�����â�zk�-#�=Xw}{PF��x�Ez���1���GQ�5���|r��4�����
��[A��R$��@m�#Ƹ9�[��0�z���U9�52���?�cG�x���<d��w����[�O�w�+UB�B�,l�{�"�P��TiD	-�3��q�h�@Z��h ��2V��j #������AF�G�_Ҩi�rm5PfŲ�*	�?J;O�aA��Q��Ո�Ǟ����SPL����܈�jh�rw�mmDz�`ޢ����z9�DJ�&���N|投���rDۂ.�<�`�d�ݮ�$�Z8���Q�+�A�D�٪cg��o��M�_?���/�%��N��%uV����=�AO*�g��+N����Ӎ��d4�O��s�SوBP~��׀V���|�֌��x��!��6Y�n=D*ά/JX��/���zV�ܢ�d�n�Y�����H[ �.�c}3�?t�O.�_�((�%ql�"�O���6ʌ�h��l�)�6.��r�{������N�@��r���Y'��G]�D_��ҫ7Ե���]�Tg������^��T?H!/n�\.D�ѿ(�gݻ�^";)+���r�:����� �����!b蒔��.H��l�M�=N5i�'�K�n�жfY��F��T�)�ָzC�)&��u^	E�^�bnI�pׂa��q��u���s)�z���XX�̨�x�4 �+��3OE���������5�P�<�(Є�֫�|]�i�O
�)���� J�[��^�i�JCo�t�?�ڐ�A�]���xB�ǉ�����O�E8�1~J���d�M��O�i�O��84�����B�wa&�ײM�ATB#Lc��h+&o��7ru�>@�f(�㷶�J�R��G-GӪ(���5�TD�٣,�X��V$�XH����}UGN
T���y%2��uM��m��9�4jَ�K�(Q�7-5�ꂭ����H6~x͂���3��h8&Ҹk��	@�2�9c6��L��������}��͌I���L��S4p@ �OT)�l?fNc����̣���ŀ>���q�}��2�o��JZ���[��x��l����������qm���]��nha�X�5���v� �\���N�p�<���-caƍ����a϶^���	wKD\^<��x�h���q�>�C��m.~˚Г�YH8���C�W|��ȡ�#_Ys��
����F����|q��x0������u���f�&brc�R��7,RLc$���9X�ӿy>ƌĜ5�3�����7<�p�P����_� �PD�A��M����fP<�X��@/����R�h�1�&� �my� $eD��R��x�kf�]���@ ����������!��Z��ܠ|�.�'6� �P�b�/�K-�ץ�=G�2�ğ �9/#��,���t���#gr�NM����������ž�5�G��CgX����\��1Q�k7I��dRO g< S[�,ƿ�^q��/}�do�Pg��d���Y�)r�fX]�ؐҜ���>W^&����-�pɂxU�&�y����7�zO��?��e��L�!M��nH,Hں�t}[��w<��b*����2s�Ӓ�l��0���p�+�͛�w��	�(H��>��,�gP�BHRKgSR�ö2���aCK�\�#.����˜�ެ��M�^�T)ٹp�n̔P��P^����*���!O���1���H�5A�k���jr	�&$�$�v�t˂Z���6x�Q���Q쥀��[g�6�l���T�%��e�I��N3�c�z����Xo�$�q}����0�/�<�9 ���&я"�����1��ߏ[�6�6�Lk­�)�y��i���6��bc&)A�sa�B$"���T����3?~P"�����w������%N[R�Jс��Y��W�/&>��GC��z�t� n��_e����u����,T��G��O%��}��&��y؈E��P�N9�}���c�j���1c5w��n�TT�UH~%�!X���V"�jI�wL�	�2�'$|����0�r� �b�0�ɉn�n�z�n������=�^��k*8��j��V2���>��x	����������u�@!d!��򌰃��ZS����p�}wX����������s:D���j��ȴ�1|��jY�P孢.��!e��C䒖{(G
�pu�?�	�ָ��xA���H����Ƭ,��i:�~���/�ܱ�܄S�:u��I.�PvX~�MQ�y���ez�RfCZL ΍ƜT9����P����a��3B����\n7ܾfVB��՗���x�&�NY5;O#{*_��tlސuP�{.҉G�%�_W>ǉt�;��>�3���m�.0;=DPJ?������Y�E�MV��Ư%�!?c��\<��?��(������f�d>		D���M�~n��\�v�@kZ���l�қἺ��������T�3'CI��2pa�	j�%��2T0�;7��7��OgRpUjw���yk��~�#b�E��ˊ���HaA���Q������k��r�zۓӬ��r�ac&�F�}�1.���tS�*Vù5q_�Z�%5U�ubi&��L�;F��\HID��1��wIj�ԩ����5�c�%�\0�����u�L�'� z��aǄ�|EU�Ȓ�=˖�Uy8����2�-A��ng��`l�_FY��N��ϸyC��%4V����g�,��+���1��Hw�ϯ\������N��W��>%��R�q��G5�S��e���liv�|~L+�i�|�ڭp軅.�E����
��4c,���}��;7��̔����{����=��:��q�I*���G7c.�l���'�T���nKFt�rb.h��]�:%����+~Q��RXň�!��8ĩ�Dj��^!'�B�FOrRӸ�(���kʨ	����x-���~�z���W�-��Q�e
@{8�H3��������j%�
a��{�S#e���ܔ�~�xn�u�Jo�ge���|nA�du!��4 1����'V��S��<� �.����f��}!������zY-�5�5�������8�`�_�_0��3+cbʹ�"�'">1S���'6K@*��mp��5%-��JY�r��4�>�B�`_y#�Y����\��B2���S~���`��Y�o��+�68dnH2Mf�b~j�OQ�[ܞ�`�x���,�"�`��#]~�hC����'�� d�(ϫ��2yz.ME�n�RS-��|��YO��8ě�;mec�x���W���-�N����pq��ě��KR%@����l{��eFl��(��-�ه�����S^���!�R�����]��ӆ6�-k1�՟���ot�VN�������Qv�>��q �����~l���r�ד�E*�Y	0	�������G���v�NB�|ogK�G�Wź�G�%�-�q�2��hTGd�$����D�|4!�5(pu��8�Q����P��i�c(qCaX>��6g�0fl>���$�Db�HL���e��ך�+x�`c
��#�l�]!{[*�5�� .�+�E�aK���J�@�#���J�B�E�@�����9 �o�^����n�gۨ���D��ߌ���m�����v��A�1��Գw旗CT�ni�8���d��	<�� �^M������Z;���hTm���{<�n���#G�tG8Ĭ��t�Qsڢ�>{�:ֈ�$���/����`�VG�2X�N:�̸��]MI��U�%�6e�aw�]�z?б�$�i�4�q7B�2��-�D�����fBJ�Ǉs�������waHv�L�0����mu�^�4�n/b��1|�i��6�j�և��t}g�|���̞��h���1s�`5��� p�F����<�3��(�W^]Y�A�B�
�'l��z��g���6��г�o�AF�ovJ	����h����V4�c��=UuL��3#� �U�gh�e��9�/�NUR��N(���6��������<VH��{&Jz��#*�פ���eC+�LS0w�\��JV�Ջ?���z�DƸ�P�9Ο�Y������^l]_�@c����8Ӱz
�{2����m�ZB�� �RuGU(�DI��}��rSC~���ݽb:�!(���08,_i���g ��E��p�V%����	�=�JV�, "�:/ ����뭑V�����偽�vc��K!�zŰ�kE�A�ZZ�
�wӨ`N�Y]�;���c���ˬ��?riG?��a����)h�-���w�4)��C��7TZ�3�����+%6������S�E��r��S�Sv�ו��
ظ�fT�dL��@:���q@JL3@�_��|Қ�<<C���!�Npn��!����_^ 4H'�gs�0<J�k3�sqWMH
I�� T�]���P+�D��to�B3"U ���wz��&Z��R�29�dHu��xQ�ꙙ���6�r8?)�|�9�|yvf�L1e(ФFH��NY陼j��3�nX2�vx`�1�[���<�e����r�7k6�E��!۪\z�8���%zb�ܓ�� ^1��6Ѫ1,0{��#�5ޝ��~�юX�
G�,���/�~g�Jd��Y��	�%Ц/'ӯ޽� ϟ��c���rc"0$��&w�v�|d���TEV2u8mz=���K������
m	6�0Յn�a��7�l�R�Y~�H9�m��܂�.jA�Q`Dg�z�E�iL��N%0�T$���]�s)�|EUz�3g�K��)ȥ��%[Q���r-\l��ǚ�:�A�X�!��o��G�P���c�O�_��C��H$�zK���!�YjQn�'��H�W��iVl- �ҾjT�2�0��P�*��Xƥ�؋������d���%�D����i}�H��}���n�S��m3k:��lBɕ����j�����_�;bˆ8��$�J��?Z��,u&���z2D�^�mgJ�ҡ��0�Y�ne,4-��M�RJ�(>] )��V�©|Q�k�-�5�TtP�t�^�$��]�I��>u��M���7�Sp�2S�8��#&jToÕ����J�It��G�+�cj�l�t)8���	�bNXӄ������v�\F�5I`o�������`�?���O|�41�����DN���h�*��ƺt��$n�O��q�W$����0uZ^����_M�1�	�|aP��oQP:g�U�����w�����4s _H�Ր/u5g�c�A�3�r�ڤnO��/�T�^���FB�K4�+<?���0=
�p�! �ڒ'T1{��������&HA�K�߀ƙ.X��/x�^�J���V/��h�3�C�$ ����ń�!�=|x�F��.}�1��f��u�l��󰲾%�pf"�����1���^�Oʿ�?6e��0�N$�Q�jD�I���@|\1@7F�vV���g/�7�����[D�@�x�.��ܜ�}TԎ��Ɖ�'Ja
F_{=�@�Pӝ
�����)Ƃ�
�,�6T��[������HL\3ᮣ����wTP	#�.���G/�9�NaV?jl�@��^y�����*����O�,��hQ�X� �h ��͌r�A=�o��^r'�b+{UO9����w�s�i	sN��רpx�pS����42��v�xg��E����klZI>%����0����d�װ`����`;�o��c�ފ�;���	��\�FDY&s0ʓN�y���-z�kц:�˃��#Q���Xaȯ,�N�RǍr����خqQ���d-�K�Xe�D���+O�*���b���f� �I� 1�I���A�RѣcןIG4 ��ٙk��1�q��p`�?��u"�E��"Y��LLeЄ;�;�b'��[G�F��]�W�el��E����=|���6޶�Y�~�u�Oz���Ͱ֐�[�%^����"��9LK�����~wVZ$��DUjs������ha{�J�����'���2O����ac�U�d]����p(0��_�5� �Vj�����Qs�	���Y���)"� ��T�
|����txK`����6�N��lC3 y�� y���U��k��4�������^qN6o	,�N&��u�ǹ���p��&˃�`��L�ʗ�oA�|�M��̭���w%
���8�ۣ��f�FQl��f��t �u,2����ٌ�B�d2�ǨͿ s�Q�|j���R���(���	�XZ�������?�o��?;RM��� n��c*��n!��D�̄nb3�V+��H��?�H���B&b�_q?�	&X�$3d��ɒ~�H&W��ç�;�<�,��I��ļ��N��$���˔X{�?���C��|�2V(���!�IM�c0M?q�Q"~U�����[��.���!�B�"�������Ss$�Լ�P(b.5L�@����t6jN(Q��NQ�ׄ_��%�6ҷ�:�Κ����	���q"T7o����0ܗ�ta�͉w��d�4891�L�g� �k�F����ًn�#�)�Ӫ�Ǹi�r�0�HC0����%�b&P�,xn�c0�B���l�"�*p���ʚA�N����Ep��=�`�z�����_,��F�sX<y��O�"�C�eǛ%��|O�!�kJ 䒾�����Kx�P	���=�}	Z�*@�΅���k�׋�yK{ꐧa��w�Θ���0͓�i�����[Ɓ�C~m`��W:_x����u�;cќN[�A\D�z19��)�@�W	o�2t»�����D] ��!�Rֲ1ɮ�z��F:K1������iS|y�*��;P�8��*.g@v&r"`0,������u/$l����,~jL37���R�aM2;;���������J�NK?�l�n�u��)�}��d��哱y�d�P�=��~Y�~�r�.0�*<$�	�PU?%���D��1?��p(I�ٶ����%�B����@��1Ϝ����kA�E/���i�rga8_����&v cǄ/�b�/#��]���y�I�C\`9KuG*�@��������t�@��Odz�A���d���4E>d�3��JJ� &�[�,�`�~��)7����jxc]#���A�'mk�7Jˣ%�C*��@����^�v �Z�خ-�%쏾����fT�3�8��SЦm*p�ǀW�`����7k�������\��q��`�6�"�Y��[��e�-�1�R�_�	�Cf�4��}�=�U� )�5�7:�)���W�fg�����9��ђ�ǌ��?`&����ƅQ�t�G2�[�a)O떳xF]�W�mS d_*��m\-�ף���<��\i�6���Lcu>c�WАT����H��\s�Pd����m��3D8.�4~�Ґu����ʴ����-W������t���k���O-��!jol�ϗf�S�syI|Y���K���yJ�0�9^�,��-f�	�Ņ�]O0�ʽ�+Y����,}6��x���F�����q�)Y~�P��{I׺=o0����;�k��o�U*v�E�J�b4�8�1'����П	1I���r��D��LC�*ks�Np��%�o���oN~�q�X�Ǉ;}gh����B~��z@ڝ�D߬���&�*��a��ـ�#JF�s��no��-;¬�A��\�qvl�n��y7�
��"F�D9h�8�/8߬$�i�9�6�y���Ѱ�!�,S��9#�l}$��F�gBf�_A�QF\2~�rFt�wj�������7��f�2�;	��P���wE�b�4G�����R��JJ�ݍ ?Wz��{�5������'���L���� �� ��
���fTQc{�|խc����1*��q�54�0rHV�S�g��I�+�J�����d�kT�t�A��w[�4}-K��)��JX�+yDq��H�`qmo��5aj�6{�D/�Rx�X��A�+��k֟a����C��7����#14�lĘi��t�,%.Hu�T��K�dT""����Q�
�<:�d��W��寚�|�a��n8^���ʥ�QM���{�����Q�u�֎q9{��1��0�� ⺧�����e������_pv-v\]`�i��m,+X�c5z�z���%�/�?,<�_��K����)����C�b9�hH4�p��.8���n>$DYѸ]"��h��=����z{^�� ֪��J�X�@�o1�S�c��O�5�Az���i�GĊ�6���~� ��m��H�Z��n�%�b@t��@D�v-_�)��.x�X�9(�����R�k�ޘ�v;!�-���͠�Pn���Yj����"�G�+��|���;�$��n�Y�{H%��/�NV�uG�&o{?m�׹k��CRJ�����V,/�l��.YQ�6����U�*o銫aMO4=6�ztN�,M[�MK��/�e��a]��ރ�Bm�$'ކ��=�.,yF0�i�l�A�B����D���v�Z.�R�N�X�?��G�8\�(���))m�Ȟ��\SY�&[��f�=X"39��OgS֤��T�^�weOwq�ĭc��R�(G-	���#6��Xu����Xx2����S��P��ˮ.�WY1��.O��	����������"o��/n����,��I*�uUa����뗧<��z���[�UaK!����p^c�X LFݞm̕�B�F8���M��J�-�a햶�7��z=��b�]�}h�`�Ĉq���J1'£���$ �sDSk��������7fLX�b����C+�����ϰ:�r�q��"�/��$���:r͜��N7�����^!���Cd~p�r��5� z+%�H��� nt���p|�p�`.`J���*����C��ᶪ\V�_��Ͳ������wm��b�,��X'��b�zEC1ׅ����^ �:ll-X��J�f>���^�(j$��
��wv�})x�f����]-�e�����
 H� )��"��j���m�;ۭ�x�p�T��U���cP�B�B!����@wɸ��92�8~M��

�xj�Zݛdî|x�����3Q���8f4OĔ����%{��K/t�O�=kh��~�����+j�v�?�+�[9H8P�վ��EѨ5QH�=rXz�F��'+`�0<����͓Q�Ks���H��7[�ϙ�]Z,�v�M��lV��௯���dq����w?E�����S��9�ك}�Ts��O!b�0�f�%u3��@l@��Tn��X	j��X��v�/l�?|�4�*f��b�d�WK�q|�AH:డl[��u$�L�� b:c�3�|���<�|�aГ.��$��&�Sr�R�D�p7�F��*�{w. ��h<	���;�'�����í:��8"y�h����16�u��O8W�[���ނV#���%��p��q�ms����n&�v��e��ʩP72�_�n񯜔��(F$$�� mI�J��pT���6��b��]�k���nT�7G�/���9
Be�?�o�����ˈ˙�}~*d	8_,��`'4(���]�'�����b��ؚ�bN�����6�A�����n�6!��g�u�>��C}#e
g�c�qV������)P��������H:�~D,`���'�ۗ�aL�?��7^۸�sp2���0�D;���ډ���=��X�������<{�e�(%S�$3����Ҭ�
�Hy��;�`"�HZ��Z�wNO��DT�U��#kZF�r��1�3f�>�Ґ0'�2�HE���A��t�p���J@�d&$��5�{E�Pf���%Kx*H�|7n��2��*����ʋ/K��so���-�Ir>J�A"�0ބi�£�8ŐX� �"���o��:�p���e
!�����R0�����f,'�p�=�h�ג���]݀�O���6,4�3F�(�n�vCO�Fo��P��&XJL޹�R�³��s�jv��%�ȵ�צ�ɦw���2~EN�] �5
��;"��_!b�>�2�Q�5 �ʲ~b�;K��sq���m]�U�{);���k�Y�Im65Hf��nY\*���K*|JA��l.�&؂ nF�����I>0m8�my"��	���-��	�)�������г�|(�מ�ه�B�74.���m/r�q"���㧡C�8��<G��Kv��^9������k��I	�B������N��bd'W���I�W�>�5�5�&�U7��S_��e��X�t��G�u����NzUÉ�5��>�@�� �sZ^4��7�����\�?5��I\��u��2����6���t��3,��Ź�+�t��X�������������A���.5Ӡc�@�kt��c��9^8�����5�oW!/_�����&��CNm�,L'=S���8�\囡'�/�f�IN�ڕ���T&���|���^��Y�l��Qj��U�PdUyl�֓A/� ���fЙ�Lvor��>�|��l�V�Rs&����B������9�wl�-+%����K+��{|Sq�}���G����;P��^XZ*U���y�)a��]�B��bw����,8s9���>�1�g�5C����(��N �a�! BL��J����(�ф���[nm�M}3����� u֌�)�P@��%�aӁ|%ΑZ����h��%^ŀ*���������O����I*�~��'���'��`@g�l* }�i�$#���G�C6 l�$d	O��J�����q�d_���	mmm�	B�b,cH�"�Y�-�0V�����0�
1�+�(e��'�fJjS؈W�<���/�vCNTuz�����,�Y{���cQG�Xv�UA�JO���o� C���%�]��Ͽ�%˝��s�i�n���.
8V��9w��~�T|6��6"��?ԭ��6V����͚p���N��F)�fȦu�����D���7�2��K�\s��TP=�^���px՝�� �â�dh
�
�[�z�N!:���*G��6��{���C��l���5��P���k�g�L�(N��B���s�t�XO8$��C;v��ݑW�ۯP3M�,��ugD��s�HRoi�r2U�V��������9g[��c&o��l�%������}�y�WO��W���\�	��Ǩ����K�$�1�<�
�Q9�)�������u�	Ep�*�8 �Oy���l�\����c���sT��mk�{=��2&/:�t-��>���Y	<Y�
�֔������,���,v�Ķq��R�(C>90D� �y,<��"��;���c�<-46���	��I��%oJ�`�*��F�i}�:�� 5I���~��,�fp�{A�u4��B7/��v&��N�"�Ši݂��&�����2���MVH f�I��{�3�M"�V"�Q�}���� R��Ȕ�c6����EIU�Z�;L."���N\t��~m��غ�:9�GY��H��)�u��0ڀ���m�-����J���)}P��Q�p�*e�!K��U!�G���u}X���}i�UJ)���/�4G�پ�%5Bj!���{!��!I��A��A!_#0��A&0����gm�����1��a��!t�QW	\��O��b+VD��49p�[��eʘ��#�U$�d^�Sö�ű��� q���W���ğ����ӫk��H�B.m!��{}��Z�H��Ğ������8�1и�ڙ�TDN}�}X.�"�=�>�6]:�����mXLr�n(MA��i�L���r����˿{YK}�t�������p�U����� rJ6VϠIN�n�G���E'��_0���L�����^�޶~W"oDW˭	(^�io�Y�p��k ���V���z/�j?{0�8v�{�x�5^q0Mvy�!i��9�2��1�<�ۦ�8�m72�
�Ão�z/�n@��A���2�ޥ;�"��N �k���U>���s�Z��B�8�6�X���3X]#2�����CE쳲�<:�[W���l�b�"!��en�)����q>��*%�u���Jܨ֙X:G�����S�q���mY2�8���L�'D�Iɭn���rk���X�i��ɢ�w���>�g�~'ɞ�($3����m�Z� �=Mrȣ��*tT��7L�����kU-x/�T���>5�r��V�i�j��`=M��#�Hy]<bIvT�=x	��kݪ*;]o�2�kh)�U�vշ
��.�������@`XKw���p-�:y��y����B1"U�P�kc���l�(^�ޡm������ܹ���<{��4k��&��"O���{||�z�����G2�щ_3�eٵV]"6�pnXF�'(��9�m�"�6օOh�Z�(�s�R۔=���E�����|n��$p
�!]q��G˙�6gV����T�7(Ca\+�ت,�V	�&mM�|o1���J�N)��S�y¨I|���Ъbz�5ȑ����cCg٬'aT��/�����3�����ٓmY�pQ���g�A~�0;ȿ�U89@v&e蕧�j6U�f���Y@
9�{�J�o��9P�?�%��C�n�\���UH��ɚX=���}&m�0VJ4Y����[GUj,�N� }���ZF�!�7��d:	��'� `��R�k����rZ(�����Y�J����8>���Z�(&�K���, �Vh"�>�5�,�q4���P|������ԋ��{�ԋ�oGJ�m�,��(U>��}��7�)�_�~�4u(�K�l��"~�� ���4MU��f�J���$�T	(�o k��V`̻f~S]빦�rY��7@.\���*���	�u�^2`�g�8�?)<� �QŰ���)��ky��K��d�����X������" =<������M6�/a�Д�(B��6�HJ��(�T��{��<�o�ٵz_#o�nTP#2ؗ�UnC�ɚ��g�A��դ#�3�x�IoiA+'�^�	�t/�i�S�5��Q�J�:}]J���"�8��&2&��*��_5�zy6n���vzp�ә5㜴���vC��f(ȇ�ݟ�sU�YC�(��U��aO���,E�,�f�tK��lx�Nك�����E'����C����a�%�S�y�X��4g����K`]}i��109L:�DoJ�L,G�i�j�����ݍs>[Ulh��1��*~T��{�|Q1�?��{�q�4��0�֑m��	2�o�ޥͦ�\%H2ߜ!�e = .���a
rʁ�����)$A�m쁇��;?ى��%��9�Ʀ)%�F��C	��R��J�|ЩO�W"&V�L��m沙��bX��n�?\���=�;�O3#z_���k�z���n���ca+@ً֞��4MW��6���(��ę��;1a݌�U���ix;b���P�hgR�?*��6	]�Ǹȗ��K����c��`����+�6�٠���@���sT�DQ1H���
�B �q���t#���)'���b��P�x�C䍐|�v���19I�X�"5��X
�+u���<b�ƶ!oZ;�����i�&�Ǵ�kA��%0��Ad�t�,�o24�w�({�񶟺D�/=w��}��x"��(�虝�6���"܁U(@7���I�0�!}B+�_�M�r�p����3K���q�'��iL�y� �9n`&����/��ɳY�c��Ǆ����Bu�-��+���6R��?����.����8�VqU����/������D��:����|�s[�Z�~׎��1�^���I��wjz�B8�Y%��&$��U��m ڧ� ���@�h܃����]����[�~��Kb�?٫�!�Q���ΡD'ùiv�ws2�:��?�QB/LaSCwY �KD^lkvdw�I�(�j<�S�)����!"�#��*7dCL�Re�%����]	X�T��[m8��a��l����U+L���,:|�л��=u
�U�N8?��2���31�/HsE�j*N�M��£�R�;Y���A��n�qU�f�8�{�̤6�o"�V;���fY�t��ӥ�y�����5��2^(�Τ����X�ZCK��7}�e���A$!V���q�_�Ј�,��#�P�҈��=�M���o'���2��¸�-G߇#��$w�դ�A�x=-/��c�gF�����qEY���;�9���?�mv^W?"����d�6���eaC>�yP�v�K��V;U\w�e�ɹAH*�_a>��*/��~�+���uQ�gZ��RZE�Q����^��˓�H�'h�wOA�A�z����L�F8�tNH���<F�@n3ݼF�-����6g��&�kI@��k�qB�f��c��9ؐr%���χB8��2�F��M��%T6@\z�i��C �'/���/��o�PC.��X�#ׯ�ǌ�%h��6�X�81ݦ�"\�-8�R���-)��*�P.@e>��(jc�4�G^7D�v?�>8��i/ra��3	�I �pr�\��Ͷ�.�^e��eC��©}Ú�|�S5t�C�=�]u��P���Zq�5@�����TZX2e���B����Y}(4`K� �|gL��ǤtT�\%��HNP�R8�!' �!ZAƑ��n�@Sh-;S�<�v(b1���1`%�����v���6Z��6�?U�u
2`Sa�+���XG��C��U�֖�5`��_`O^s��ey����A�ݘaø�.�Px �	#p�v|��;8X����쟶P0������ ��2�:H�+�(�`Ii/8��.ߤA\�3q'�k�xI�】���u�8��֖��|T�N��B�5P��wO�p��yq��S�B���z���3g"+e�~詅p�+�\x ZfA��jm�6윆��n��;�#4"�C�C"[�WA�>p��\�j�\^ua�q��$��I�S�y��m�t<&K�^M��"ݚVf�@2)B�M�؍����7���F�D�p��n�|B�����ߡ������	���P���v��x\Z49Z`6�#���xGZ<���)��Le�k�Iy"p�9��٠;���fKw��t'P��xes-���F$�(�"�v����^�߯'���2���%�����V-���I��}p(��QR�+�;/^D;C� �Rl��6{�E�r�Q�:��nGQ��չk��J(��>M�����һ�0�K'�Nl�3l��,`֥�:`���������F�C~Ek�j�"6�`���k�|������}JIf@�?<P%W)>g�#_��&�M����B������^2e`�U�y.ʅЋ鬀q��@��1U�s�����a�4D�ؗ=��*AN[���3N}`�c�x�rnꣅ�A�C��D\8�� l���uK	���>+4�y�r�т����Or�aI�,���,-ǋ� ��a���ђM�<��ˡ��Y����]�.�x�Hb�ڰ�/�����FD -ۥ�k������5��[����Y�5�� ��y�
�-���|fN���U��w����%*%h�s.�$Լ���l'`)��R�>-pt0nib1�(�n��2]��9g�@sV�w=^�bf�@����������N�g9bmx�R�S1[�6���a'E���I?z�D��;G�IY*d��N�;��V��L4��ҥ
�@p���Ū���W��i.���u�Z" *��9Q���'53�qVL@ݰjX9@��`����B%���	C-�rs�WT|ʿ��,�\�D��ci���7?_yg��,L� �͏7���#hѲ(���=��3�W�0��*�F����E.�VPVh��u�fdr2.��v����h.���j.ߎ��qv��v���/]�Y� |�W���b��n��D�9�SLI���ئږ\�}�w.~��^� <Q�;������Op�%� "hd��b��7�U`>����H�y�����4�W6�5�e�R�xۿp���&�7.�HQ�N�"��m�N7*>#�h��!r�7'868�X�Y.hO\>�y+ld�ؠb���ēj*�xE�y4�-��cׇ`�2�9���ѫen{kҡL�A�d���%
�''���|����3
�'Rv��?���'^��8�e�����ö"��G�U6�7
�O��̑��{8�ia?��plg���>����9��1����������Ǆ�;��>�� ����פ���V�c١�{Y*� ������)�ҤEzCe3q$�^�8��t�@>��u��t�m{����ӌ{��u��`��xF����ѥ�d������f�㒆�x�n�9�� �2+�_��8��:4:�R[]r8�����ڗt��ښ �����~.�#���:Ca�?��s�&߇c��-M{[\���-p�3��E�I�XH��(�⺡Ei;�r���N[Z����N���[ �x�L�^�;Z�����p~j�Β���aZ7�!-��p	k�xP�fS��|q8]��E>H�Z��\�{W�M�=ٹ*��/��8*f��Br�����K�`���Q`wx��1K���N�%0^H�G��b��� �hnfZf��y��^ˆ��=���Av���7�w�^�CuX���F?+'�������
nV}��4�yz���7b_�A��}Kb�]'(������w]�6#%۫��Ą������Sc% 
�j7����*͚�p� l�Ff���j�Pi���C��Sc���F��b�|�8�Q1=��<�QG� )2l�V�*�J��ji�# ے-v�@PC����}�(��"��6UkP#д<E�]������-o�,��__>AI���e Ch��$׬����k�2C��L>k4�H % �e��Y�~D5�f����Ӥ­�8�Y@]���/S:r� ��ҡ��c��ꔄ�^G�H�z_��$�{=d�
n��I�6��,�����f���?e��!�<6+��c�(�m����'�	�F ����c+��E��/
��Vٿ4:��5w���7��{���K ��K)|�E��X���
������ن�30Z0�-E��Uʤ���hQ�t��J�{Fv���sbK����&�zh�<~}(��ܑ�,�T TՕ�Km�w�F�=����w0�E�VAƒ2��S�� g�	v����Y*��|$��{�.y1�P���n}��ŉf�~�H�Ԝ�	y�Ҥ����,����q4�.t���a��9��.7������N�R1���h!.һ���& ���+P�ZH�'[)dQ L��e���ſ�f�=�}y~w>�c$��v��+[�>�aZ��"jU=@���릋�a��6`�K���&+�u�廘���8$�zg6_/�oO���!O�V�/�r�`
�*��H3#�%�eP��|�^��e���+
R誋P�|1ٴ0��k���\���a���:Zh�@�B�6��	�g���BM��ek8Y@%�jW5����X�>G�K���S�}wD��׎��P��#���!���UYR�� ��'c�r���	a�feT���\I}b@?h�I<�:��ʑ�הo�ֵ:-�[�j�� ��?��Pn���?�e�T2`���C�:�&��9�x�&!�0���7��4/�����y���'��2�����3=��f�Ga����Ƀ�{�B綮��"�ۃ��s ;k���S�h�'��~'�ȕᏝ�ё^�HGX�fS��g���!�L[�����F�s��n̸���bԟ8 ʘ��g	Ŀ|�Th�t�2�N�/>v��\�������U�R@�+��l{9�o��@,�6G�*U������f�÷A]7����M��g⏦�A�_��v3��������a�u<D�k'r�y:�6��>5oڠa�w�Z:^p�Lh�*����,ń-��}��_���+C�1�o�0�&1���T�L�_��|����@d��ߊ��8`�u�y���X.x5L'��q�2

�-�K엫��G���,�'��T�ay�t�/É�*8����<���&y1V�[��բN��SG�FА���7f�*X���--�7,������Y��e7<�b�Î�-M"�MS����q��볞��תS+�R�(�]�;V��0�O��.�o���f��g���푣?)���9�	�����
��N�M�u^�	�Sݮ�_gG'�����7IzC�����i��~;�H'%qe�6|/��abtB �.�7���)��g�B�r��`���o��*قa<�<�wp�ݡE��A����%]I��Dc-<����PO搒�a\M�r'�e�.��㰹5NG�QC�Dk���!���is3&�0����䞒���\������ĺ�����4�<�b8b�j�EtC�(w�S"�BmV��˹:=\æ�3�,�2o��^�J{]�D����r��m��P����'�r��>�����{���48c10;6�f���4>)W��M��Mv�D�[i��1�RXb��$�m\�e�'�\���6�;	� uF�)��|fL���0���w���Fg��Pw]5F���)�F��������V�fg	���3�m��CZ�l����=� �L�qYjf�{F`

��D��dS�JS��R��^U<��զ��������7�|���Rդí��%j��b�L48���]G��I��ɋ�`o���q�& �Q�m�Z)�G�RZ"�C�̿~�Y3���U%mKǝ��-g��}����2�b���
�2���n�����~����T�毭���p:~��RA"�ķ��{0�W	Vr[�3+h�Hr�p����	��e�-�*�ǭj�GS�':���3C�D��A�'|��(+)_�!����!0�Wʆ����##�c�m�"�.��
���x�p�1���V��4�(��nPi	�����
��!Uj�.O�ix�
-p���D��GM�ؓ\��&Μa>s�˼)
��Y���or�>��gW�*'��L��w��j�v�E����sl�2X?���7�O����q5���b����u�m��4�����;�x>;4��W�c��ʡb���NW��<�^
�jFI٘d��y���&,�*[u�Y��/�[���L��ه��#^��J'���ޡl�0���{��=l֭�}T�6��|p����{��
�!�������PN�}bYD���b���-��d��[��˫�B�N�sl��C�f,Jc�>(�$
&����;o�V�ڠ�(UdŐ�+G�98-�i�cҖOԞ�no����4>��4,��Y��ĉO�)��ka/7�m�b]��7_E%c�Kx��]v6�@\���ᚺ��:�������,a�g��b<��+�[c��|�sȋ���FE�3��j��k���@�����F �[*���*�Pf�1��4���s�;��_�.3�bl��К.�����Oڄ��g�a8INɣ�������?�b�JZh\9YlxM�=/BVĔ��h(��f&�Ү}�L-�{�ɐX��D����U^?�a	Բȱ}M��o��z�e�"L���ﾉH��^s��YDy�ӣ��j�MtG�xf$���J8�[��|��(0���|;RVt ��<6G�e8��>Y�Ҙ>�I���$��3Z{ ��
�]%���Mmh���R�>��bN<5q&��vK���;��	���F��4�����i��c(�����鴦 o�1�w8c�;,������?��o;�-G�)�h	��m�1��.�"��2������z��ض/��ɼ9�	R�"��S�	L`P�㰟���#{J�_;	]?ۊl]ҕU�u���>7M�?�PE���Ay�3~��pE�m�ش ��
p�o��9e<�q�l�Z�,i塵*Ҫ�Y��H't��J��ۖ�P5�w��o��I��9o?���wV��a�9�3DEjŴ^S�ӨI�$3l+���Y�(�|hg��+%�b��C�EJ���!%�v��w�6�pYj�EQ��xzU�*��\�H
g*���
�kc���W��/s ��u����,2F������/�A��Z��x�*�ca2�5���-�˝X�b��?�W�X�)�9Q��8�<H����r�X^�o��쩭J��2摕br��@��-�:o*�iZ�U�{0Y2s�E0~�p��AD.�Aa�n�SM#m�@qՑ�^�>������ô%�Ѐ��+��+hCA���+x,,ǬW����o�6�@�۴҂I�"�~G��z���c�h�ab��J�/���Y�D������'Ԉ�V�7�3��ig�2���X�_#_�"���>RQ�q���5�\Ł�V�j	�l[����޸��6&aZ�%C/�z�!�GE��*��cG�d��(����n��z*����p�*w���f�	��x�O}�=R�����+���Jy��`�ID��:� 3���3gx�Fj}`�L��#���D}s�j��3WBʴ#���uIi$"�A�>�~f� ǁ`Ž�.O�𐁨Ų������C���֚�,t��z�k�$]�֞
I@�
���l�7gAu.J��^�����Lҙ0�؁�<S�����G[9���}��n"`v쳻_]<Q/'�E�nr��(�+p��_?��<�Ɩ90�6�.1oB�
�~��m��!�f'9�]���d��^Fi����GNn�eÛn��z���]�x ��N�q�c��EP�t�T�vaxQW�^�#D�Cb�� �h��h����q�OK6����,Z՝s����U^��&�"~�D��dTJsښg�wZ'��)�z�L~|��9�4�&E�+��m���^P{O)�1y���*Yf��~m`~5V�g��}�{vev,�n��e�U=�y���AX�j	�
|�7'��P�NW!�|~;�j� ٶ;x ,Ճhzȃa��'䷈=�����v��Ox��{����2�D'�{X��ъF�+u�S!�^L[�T1���1��d}�g5��OHlS���:z��4$��� $�GDo��fvv�$���{��?	� 2ai,\Q�C�,ee���#cS�<����=Qw�D���N��Y�=�~����{�ܬ᭴�y��շ�%���s1r�(rc���(�R���k��}_�ޅ��x�IZ�5�	��������~��sOXʙSqV_{�i}d�rN�1!z�m�?��F�HV� ��/�HG�C�Xʯ���	�p�ٞN͟�����3TbD��V�'2�qj	zxX@�=,���M�di!���w50�:(��B�*Q��gh��&�A�!�Z��V�P�4#`�~e��˲+���Z��V���6��X�W��ZY�����`oF��94�="ى�P���{M<��q��n�O>r���7ȶ�0jT+@��ҝ�s�Ȥ��h���� L1���x/nt'mO�1�1�B+J%1�:*<7���xL�nvͬ��1'�ٗT@:&&�0�L}�;�"(T7��ŵ�u�(ym�ǋyH�ʹ��(��5{���!���_	�;Ԃ�2�8 F� ,���W{#�Vl�r�#%I��F�h3p�K�Ӟ�m}֨
g��,��|˵t��)|�|S�ݜ�Z{���t��uES�Z�Aq���u7{��6A�G����{C5��Ԉx�ǁ0�e�i��bV��������� �Fn����z��-���sv��|# =�zĠ��,}�,�Xf���%[���T���a��>�\���� ����JP�`'H��̛�&�2����ip��-_�hҶ�$WxA���۰`����x۳&R��:�Bd�����}�6$�>��dH��Q �b�L
��ը�*��M8��{*�-Qm���lhL��}�3+R�%2/�nڇ�3�).� [�\lo�h��.�ت�ij)8;�,�����So_Xȹ�U��r[D�9���@�
BD%���_��7���v۴�(X�[��a�T��膉���?'dt����8pzE�}��ڭ��FL����kOr�۞���m2Ϙ��5��o���U|a�Y�Zd�M<�*|��	��+�nf!��v<7����[-�d����������9�e<�@h�GѴ3��Ąj������S�p��4�N���\;q�7CW�o'�A$aL2_����H��5Yw`�[P1,���HP?
`3���|��MMDB�ӹ�.ξ�K�R9�Ik���BE�HP��P��f�V���7����x�`�aV�D�-�C�9�az��RҨ�ڦv3�B��{y&�/nD|���W9��_:��K$r"g�_ĕr`�n��zje���}���|��i��gU_���1{��b�Z���1��,H�����U!+��R�����)f.2rB_�?�>�&��QH��y4yh�j���@���g�D�ڻ�<|p��2n���P�eJO.��%t}�P~c��{F�Y��yaC����x�1E��3jv���ՊM ��Ʊ���6@��sS�-�i���?|��u�q��8v*QN�e:'�b��<+rF��ɞz`��C�5��K�
������<��"T�W=t/���GY4�_Jx�r�~���ʨ�����_�[ې�z5���N�����s�B�����CHo.">�}�Gp�2�$e�� �_��`	�u�a�7�t����.�� ���)	�q�=��ŬvOYQ��P�f���-��ͱ�`e�*ذ�_���Ï]j1H�'��T���\�r!��ʬ�r2G��
vH9�&��V��k�s�i��V��K�|K��o2��:��uU 0$X�ۋ��_sb�K���(cl�q�L�]���IӸƀm响`�%o�_VUp���3k�����L�V,�5�����F�b�}i�0��Hzmљ�d�e�=�ŞR�x ���B#�9�g`@Ỳ�g2�&��'{�@z��� ud�c̴s��<�K}�y;���
�޷7V�=s�6֛A���Q�6�$x⬋d��Kx[E_�e{��<�&���%`b���&�\�ޝy�J�I麹�N���M�Q�5�h޶�!�J�?��8I�\|>Х��%}Yē��26a�2ُ� U������R�E����@���D	�_��@���ZC,*08[�՚�tAw���J���}'�6�C�Ro>��E�u����c���`ZC+ve�a6����� ��󂪤C)Kڱ��8�WPE����O�p@�i���w�+_fG�H�0	 �H��A4�ƣ�����wm�$��n��<tp�&�xU!�u��U1j^��D����pMj
����� :�C��xg�^�gV�@C�6e7�)I����M�mӡO�s�y��K)t]��AT�?ڍ,�==�1�P�h8��#����?3��SF��)1��f��kh�|�C�3��[�8���-���Р��[]�r"��*+�s�#g�Õ#�l�� �o(�J�q}ш�x}o<q��1^��i}�夝L�/ͪ,}נIlGpV��=����+��F���$�� �@�r@�x"�4d��	d�JX�t��"�6�:B�aE'�b�7.��4�1B�ޏ8v����0�L��0z��=q��$�dԾ�!T�G�����m!!]��&��>��_ <ך�?�b-�b�/g��IaА��cM���V�����V����Ij�_Zk�
��ᙻ��3�N��I�g��gS���8]����RkR\��u��Сm������,��~���+T�5�udw^�9vU�#3����9��:V׌����V��NbsRH�p�)�����B�y����j�S���4(��S���ðNυ��R�*H�RY��$�zBO�U���1����_�B-�?��B6�_ߍ>��Z�HQi���������H���8���V����јvaaU��scZŐMV ��^J5��j}ƿr�(��Fi@⻳8	"`�T��UQ��>:bb�H�u�	�Q��u¬�~�K�m"�{-X�ܫ��+��ٝ��l�o�b%N��U����<sڄHp2q��A"H��H:���C�ބ���F���E���� vL	Ł�i������%N`�,��E��<�DY�pWQ ��@��g�ꎗ:��䙩+�μM�[ L�0,.�WM�a)��8��R��9.����sx\�	������<Z�ܜ,)�]�GČ�T���TO&}��sd�a��j9|�Tb��G�z�a@{�d�C�*)v�nF���P&�1�?n��g�eN�f�� H��vy����r�c'ju, ��9�,�d��ޒ_>��h�F�<,bװb���U۫���;��J)'nŜ9C2r�~ԝ�^�;���ݐ��z���?��.����1� �[�z{��$F,i�+xa��P��t7�D��h����JHѳ �[���m*~��ӊ|�0��=����0�e�٬΅z���d�h6]S��(��Ԏ�|��@�B`Ju9�Tk#�{�ɕ�"\{�u�>�� k�P�~Uf�kYCD�u~����<�Dg�n9\���0�By���?m̵7�����83��G���.���������F�#}>�6pWf�̨>*41����
C�U�ّ4%������虘�j.4��f���]|���0t:��Ey�t�˕�~M��m�g�w�1yo�_��o����a�b��ņ�t�-����.����
��5L�B[��f`���s��qU�]�ti��sʆ'di���F�Z �Nv\>�/Ѻ(�{uځ�x��y�E"����	��E�,�����n��ʴ��i��[�j9�5j�k���:'�h�j�vۤ�!W�`�ă��{��ד�M�gۡ��JkH(05C��p�YU����0�K�t ��������ۿ��7�pG����{����+��$���0�X��b`�K�����2w����v7(F���XRK��?c�P��R�U`���6Z�g�qĮ�`����;(��e����W���C��sxB��mQ�#K�x��h6��6|�Ϩ`�^�3p��=RWC��v�v~X���J�cf.�f텊��ю�p��@������;T�F�L��3
M;�j��ӷ�Ăe��-�~Z�vџ��Ը�c>�;SR[3/8O���e�xMƜ3`e?x(�>=<! �-�rF�F��r<<��</�مiXY�.��UM5��[[}�Ǌ��=�v����F��$A���t_�X�ߒ8Ustn�N�{����®�M����&iMʒ�d5�Sjc���T�j%e/�]�����#���_b�'氆�B���e�g G�C���A�-Q�J[�oE��* i�ȥ��|d�V��0�^O��Q�q�mh��O|w�'�V�kW�v� f�=�ge�����`���<�:���N{1�)ĳk���Y��a5S�@y�)@j����=�7iE�������}�12B�X��l>%7�Ju�Z�=��䂙0F���H�O�Ɣ���x[eE&���J`x �� 11�XSkP�}937:�D8nԧ�������hOw�e%k� �_�-�41����Ƨ��Y171�$���MR�h��梶?��!� .hi�<�1�pT2iP�Z�8n蒨�<k�����مdk"2�O$��5"�P&̲�U���y�j�^����;]��z�S� ��r�R
��9N����/��U����jOfק;t
:~�b�2(��_��w ����9HN=kfo��>�Oz�n��L�_���X���&Q=����@Y�R��8�*�I�5y@��dZ�oc�{��Kl��!����ΧjF;@�^����n�jA�N����Z����]�C)U�>�3� �M�|ѫ�cZ3�0&K]V�	MCX#��|��
r�3l'��}������ls���(x�]8�0j�Z�ڔ y��	:m�떻� +�}b��H@2��߰��:y"�te(�`b��9����_k_��x1����<��u_����H����5r|��z��ǫy�V���Z���Y�2d�bF�=��x�:r�����wp�tVzW��nJ���8�{�<Eٝw�1��8:�~{7x�2�+(���~n�DR�k�|��v�a!����W��θ�*�l���5����ClQlt������5�'���I��YE���������?=�T>ǝ9�]N��S-c���qax��w��ㆾ_�jU3ooҭ?�j�<��*v*؞z��e�Y)���5��Ԋ\}�n_��q[�C<�I�����ں	'D������F��XZ�bIծ;���>���Z,ա�|�{��FԱ\n광66�o�%U��f����?P�?$�2~
�|IXN@d5��h�J��*�=��F�����0�U(k%�]���
�D%ar�&��M�ό�N��
�9��)k>�mH�k{�W$c0 ��ڑ�ݟht�'���)��_"]So��Hc�3Y�ZDm�<��D��{�C�|��^ ��k�!-��UW�+	���`�݃0k����q���*�G�꣭O�Kh��De�BUBCoa�"�����]~~��ل�_�]o�7�#m���~��$hʡMh��کi����m��R	�l����6kIk��5�����h��I+Xz�h\!-�˄����Jǳ�Cu���թ3���i�,���lK��*�=�o#��
x�gX���}AMY�J��Eqؙ-�%UNG�^*D.Ѵd�m�,J���1Q��j��ς5,&���l�	;�����A�Z����`��n�j���]g�=Z���]�Jhb��9��ݹ�¸@�3�T\c��9�2�I6��8���ô~�:(YwJ����ũ���V�5�Bz�dz�v���/�D�}��/>YF�+'M��y�ȟ�"F�}Q�����g���|�,�oN�֢�|~:3���f��I�Z�5I6f�ZBz�XI��G�Y�����:q�M��O9�7��m�٫8�L��C�~~a����'(��������L���)���6T϶	>�(HC�)���^#u�r�\%�5��w:�� 
ԪA�h�e�-�,n�Kqm�ѢC�����Pϲl�d�-�"(L,���G$��m1�g%B��쫿7ދ�q����n�����T4#�p�,C�<n��[��ۈ�5�i�yT�e�����L���{:��0��̣oh�R�]�5��I���~*j�Co�4o��#�F}��zo}�k�� X���Q-�eN9�w����k�	��w��F��f��ak���H렽g6�De���
/C y�M����%Y��<~\��K���S�Z���
U��y�9�⟓nV߷2����T �4���.m���D�h��RKRF��W�?R�;�*�:7��`
��"��uUC�?�U}S	��MT�薜b��jri�����{��衕�d��1:��שC�ț�ھ �ٸl�?�o��n�s0Wh����wO�MK�c�}ߔ��k��x,i-Vj�o1z/�Jf����o�F���%�6�\JQ���菬�����8�dvn-9($�B��'���'�z�n�
ݯ���U��M³���i����3�V4PP��\_5�49g߃��ζY�m��L����Wd;�NE�Y��-��`�/ ��|��u����kڬR=�����[�6e��h~�D%�t�x�G����a�x���w�I�SM�ҭ�h{3aB�M@�BK��)�����7�������[�^Q��a���[����fq��D�m��@���!=^�(�O�j�]vE0m���Փ_s+-i3�6˹T��:z$n5�<�P��󕿹w-=qZ�jV�%��v>u%�1fx�� �ܸ��}^�!\�[� ?l�J�d̹G���c�Ft���Bp����{��򩘒%��D��XeF����v$_�v��;���L���A�&��!���" >�C��IT�Ĺ�0< g.e��S���=5�{`�z/��3x�<�^lIǥf�0�~�G��);2�`�{����tھ�9́����� ���?��*���;ޝ���k��^�{�	1>��1۠C�ɡ>�7�g�5_W�bi�
@y�߫l5��e���0�;=��s�)�Z|t#�[m�]iݾ���Й�6����htR��9+9Ux!������?|~��Ma��)�/��un�JA)i�Ӊ6�ֲ�8@�d�!ڹ�WTh-pq|)_�:��S8��y�O4g�
�F�����@��ťv�r�y�gH�{'�|���)�m,s�w��vj:��P�F�Ȕ�OZ�~m��s���"���`�u�#�x��4&�m��bJ���:G��|���4�$�.���P�H��+��O@J����Ѷ��|0 �fEk�M����B�����-��%���j� I����:��n���#0[�B���u�=�֋�I�}NW'v��7u"���C,��5X���P�_�0Yw��,�+P���#��m��7�ph%�`�=��+jx�`�݀̂�x���lf �-8��o������+�B���ıi� l1'<<����M�dJ&մgWk�N�Ff0� [��|�C�dM6q7�*Ia�O�6)��c�Y��O���w�p[�3odL���5Z��w�v��v����3|!�yW����H�� y�Q��
G�V������wOf�6Z�}O�C\��O��Km0EsN.h2�N
 ί0��[ M���G��Z�8/[�M�W���&A���� ��%�I;qu|�Z���v�>�_���k�dW��.��hMps��ɘFp������]��ƸL�0um�&r�[�ۉ��!�N���>Rkpc�5�,Py?��EC-ϵb�'�?<WlF��M	�ƍ�n�'�:&���c���4ory�vkh�W���	�L�Gm�@7�E11�UT�lT�����R����P�����-_EJ�[tw�{c�`�H@*Y��ĆS@�`)�������A��ǹ
跇�_��Q�+�@�m�9Xmҟ�"}_o�<�I��pH������$�X�~'��?��%qT��K^ЇuH~��	�9�R�I9 &ug'"���c��%.C9�L&xb!$��22��ʫ��sS��
���z=��<���(��l�*>�vnY�l�y�hIr��f6|�\�����*�s_���B,a���S�-�HA�V�#p�!k��V
:���|�)�Ӽ`���\Bz>F�7RT�d*��"��ѷ9b~p	�3K�2�f�L�=^Y\>�����;����lq��5�`��a�lCņ+x��O��nK��H�)M9+�PeG5Y���~�Jmw�.�7����bbS��82 �s��m��N�ӇA� �-���;9��f4R:-žfR��āS�{��h:�H�Vh[)2��9e�P�� ��ͫIUW4��g�K}�5��
'}�V����Lu	����q,�������E4u�|�� T�s�@���ʊ�	�#hV)�]��>�Ɩ�F��OQ_1��E��	�y��f�UȔ�M�� .'��"v{���_ũ��¤�����D뀳-�a<���t��Ë*� >�J��]uE�����n���ҁ�Dc�9E�@�LF�)�Tҿ����<Ig�����qp�R-c�&�?�tǂ|�<��eɕ0J ����8��Y����*
�t*���N�l(��!e�*F3��h��U&*���4{���2r��K�gp	���Wj�a��Ըr���U�I���RM���i(^����l���1�"Cewhv0d�2���ò�+�Q��^P�h��!��<&$�7��]#�8�l�?5Q����~O3�Mp�(�	-�i�+�$��O�2�g꣑�x��MK�E�0�il�I�#*�8�PO����\�B��1���s �7�G~P˸=kG䵢�D����[|wl�:���"�k�]�
I�y4�����0� m}7���I���@�Y�ߢ��@^9���}����M~V@j�@�W�����!�E��Y)\c" v�J����ϝ�Uו���?�n�3�0U�P����"�����0��^a<&h8oGE�VK�q�3�<�C�� p��um'c�0Ap@��h����ɝ�(�JB�
���������b��2��dB6�-���b5��+&B���Ԍeh����JAH�w^¢Z�v\�@>
Tb���i��bx��ʁW�8��|�;�μ�O-�������	�?�C>���FVe���Wð����?�OWt���,��HǢ��^�89�4�����ٹ���Ys(��_f3�Ӵ���zRr�{=��)�����e#ك��)��	b)	����"���?�RQBvE��^����G�-� ��zX�<|C:#�oPT!� {����~_*��F�eQ��zy��� �F� ��3mĩ!6���d|��}#IY�8��ٮ��B����KD�x����ڣ��<��'�Zq�����W�{�0`o$��)���2 *��=��W���{�ƃ�Q�k����[��%N#�#G����H��9)�K5�|��Ҡ"��{?���ԯ����`W^O	�����sI��������1 �+j\�⌐����P�X�[W����(f.c"����Q	]O;x9%n ŘД�<���@�!�v봲�D2�nYσEi�ǜD����X�f��-�Ɏc�n��D������O�S�X0
�䛱$(Rz4��PTkht�����p�����^���W��<A��/�OE�R/��A,���/�R��&[V�0sf�N3���� Ĕ��n������ (cBt�w��:��/"��1w&�_>�N�������7;~��Rh҅
~��w#n��"q˺�΍4K�Ɲ�pڶ�1K�h�9��Q
n<w&2nKW�*�;ҧx1���I����}�zf(O��V�<Q��6r����� �Hg\d���1��Ƒ /ڶ����w��铎��Eͨ��ư1��)���e@���i$=A�0�k���J�''$�*Ww��OH,
w�i�5v�.ًb��·�L{v9Cb.���@�4I�a�V��:��FH� ��0|�c�ef>�������y;���WtMXP�V��ō�_{��RG��?M�����DRҪ1*.�ws"<a�H )��f�U�j�)�@���f],St߄�
��2�vD�im��Z&[v$��tvJ\KL�֞č#��qIDS_oI}:?�5���%����uD�/Ky���Aj+�;�>���e?҇�|���Dq눽��q��m0���Dȃ=
��wA,�m+NQ�Ĩ�0&��rk�Xi�V�m?��Y&�H ���YȭZ�-�y��W���4^�uP���k�Īi����^#gb]����x�b�q�A�Q~ZP�1(�J�da��Z0x体�c�Mv�3��� O�B�8
�	�K��z�ᄓ�a�儜L[�@$l�Ͽ�W
g��p�߮��u�� ��'���
��c�5o�A���k�6\�l�r�c��Jx\�2Ed�/S4�_n���@���~>�q]��Ӕ4,�6�� L_�Tӵ��^��5Ti���.��J��� Ӯ�#3?��uC�ܟҚ�㺡��_�.��Ij� '
���W��Wc��x㐨|T��MҠ�OУb$�"Vz���'m5R��]�zv/`�lE�K`U��b�dV·�+�@=~���s�*r����y�o�� �����,��2��Z_s.�-"ѭ'�.�0�j6��aZ���W@�@�j�F1���R�;���w��4����2C�?I`Cc�{��;'>4'�NTU��I�Ds�� A:��.3�6����Q3��	'0Jv:�FI+ D]X�H�]��u�!����0�w��6���=�)�:�ّ���O�3n��D)<}mG��Ȋ�H5G�UD���ǭh�����?�C�����p��V#&h�
鎱m��D�u��]��Lŧx��ZO� , :S�@��f�%�sM7 8�:c�!U!��/=�j�Y��Xi)d�Iwu9�D�4�;�VMS�dX,,K�>��Ĥ��{�:�#{��ɕ���R���j��Y(p�@(Cmz
�#$�{��w�' �ѯC�O���������u�լ6���_���^��w<Q��+���`�54����x��,-�?���i�F/��w�nr� '�������Q;��N��9�U/*�um����is֔wb�+i@���.�<gT4����޵d\.���;
5�0ƪ���E��l��Si�#h�>-m��2��m���
�k�i�?�$/Y]	'�d4��`J�[\���}�9¢*.�����F��`����.I4�)�gB��Qc?},"���-23�+�܄/ظo��6�~�Vd��QdS��I>���s��58g�r��Y��p���:����HyD�_h�MH'߫Dn�Ofe����@�Hn�d��y˚�_�������`���N�#A����'7�<�?FNݦZW�c�a��|$(Fv�F����L#��Is� � ɡ�m�n�U�V>,�	7X|�e��]t�g�*�5J�f;)j!�|4�[Q])����Q�~+B�W	&�`⦳~��ʨ�*���O�aAvY��<d~I�yj���d�m6������;��σ���sw2���	]cт�k6�W���Hw=T����ꥭ&���u)�9���yqZ�Ӑ@�Daa)�w�O\��/4ԛ�.W`{U�^I����;[e	��$�ƒ����K�XFC���\�r���:Y�OK3epDǫ��3Fٸ�-J��i�jaCHP��`=�֌ڮg�r�W��ǺT�l�4��zk���RJ%%�0���T2�1K-T�J~�t�+�1����F�H=9Z���L-o���.ı�B�I���T&��9��QT�,�'o�K.:��Qr���\� ��)<�Wi���%.�%�B����*����7`u�e���Kn���
�V�F�m?N�~���2㑸�i]���r��p��|u�\W�$��y�V�P�z_3����pD��D|���s0��c�S+���J�����7��_�#j�yrh�<���p�0k2�xPE�
���p@?ĕ�ܦx����L�E֐��3z��o�m��9�/޸0�QAB����:��F|vV`��̚�v%�͜ω.܌�ںo�<%<uU�U���x�J�$��x��u�k�x�ތF�A5��a��4�'���܀Ξ�i���:Q}��}�@[������R[g.�>�+�iF��R���2������<W�L�G�ml,�_k�tY-)[E7G}&A��^.͏�~s�h�y�;�	�����ss���*)���

X� S��A����zt��N_V~��R�H���.G(�"���s����d��3L(Xu����>5��`D�f2ĸ��L&��Y��JA���=�W���R���V?��q[A������y`R梤./���~	�k�ه�ب��	�\�;����Dx~�F�Ìޙ��7��>�b�a�ƻ�я����6�	Ы�A��rݚ��jT�a��h��.��||=��@+�q}�1,�_��������♼�ה<t)�w��M%a`k��j�aI�J@M��ݳ<�װتt��>��f������a�P������a!d���g��0��]� �e�Lh��W���Wn��p���\(� |E��2�}$3�؋�� ��BB���]�8�_��e�lͥ�s�.�M,S���q�ɞȾ"(��uL��dGUg+	-��g�������5�H��э���n3;~@(�H1s(�ʵ������$t5%��� _e5&z��G���&|�Qj�vQ��l�}Z����o��m S�r�}�_�����!)��-%|��
������4k{Зs ��&
�^Y
���p����b���&}���7���P���_��v��'����
������>L�k�DT��q�Q0�7XUE{H�h�^>I����}�24D�t@ڈ��	Nc�`�\?�*x`�֠hD�s�`he �O(b�L�2���n�6*,�n��M�Ҽ����2��<�Z:N��w�D(���w�j�zp�yz�Rw�~~q ��-�Vt���#����ަT�`
�R7b ���;%q��@�T틙n��mj̢��.E��0K�Td�k#��:�����b!��Ok'���1�LW�D�E�gE�h�f��D	��&ꋶ�+�6�"@l�C�f?�	^�
�Z;�$h�f́p�a�r��[��5sҐq�����٠w[��,ձ!���z���+~+���e�x�\��{�y�(��8�7�	8�����
jg��;�T�J伮�=K |X���������g����pB(vg�TŌ;���xʒ8�T-�To��dyڇu���G�F_&F���\ML����Y�)��0œ(.��n;�Cg�ŠT�֢�U��6���q]�f���gE��X�j|��R�S*B�O�i�0��9��ٺv{�	�۾0�������Phߴ����콝A��n�]$!�\-��CH�&7�嵎�@�k<��h�����*q�� �T�Pل�x���C����F�T�SbsFu9�㲔iu�n+�l5@�>c�;JL�b�P9���~A�*�
�`����F<���_��+45t��C�M�N��1���n��|��6�~��ߜ`��r�N'�&o�<�q��9�N��~�O�[�>��r=�{����I�գ���ȹAV�"��%�S�׭NT�ɋ��Uz�?�c	LV���܏"$�C�AhC��ȷo�mym}k��&�|>r����s�A�m�!t.�HV����rWA����J�W�#�x6V�����z)qkMΔ�;�ڷ�^�6�p0�b�Pld|����H����"��X4�X/�0D�F���Yt�	O?�I�T��=�R̯M�:��`�7�3�T���iB���&*��I�Ӄ[#�;W<~�u���I%�����!�)�ZSݽ8,Ғ��6�wM��ް�a�`��u.��ϸ�!a�K��j����t��L~��E�[��ċB}S��j3���R���t:Bq��]uq+Z`p�gU�YPau�#�t����eth��BQx`�H����z7��:۾�������i������o�	`ʱR�Ԙ���<B�a A�R'x��a�DG�k��H�>��i�
�su�����~Z\��\z 'w����谱�:��Q�i������fzZ@}�t�(�
��5��	��>�@�@B����UViG�UK7�� g��{���*Hԣs�{Q*crg�ُ������
z������Lm�W���id�N�����~p��!�5s�&0�葹�yޑ�]��E� ����*�=;w��-:���зs��0$=g�̥�<=�������
 c0:�dq��D*�\�>[��wİ��e7Lw
��s��Ě�j�A.��,v�L�4i�-Y� fQ�l���(u�Pd����Pn�xD2?q�q�C�X4C���9�U~�뉘U��<�&'$�����rбA?q�q�.�6!�9%�>���$��t2/a0ddhJ�me	��)2�$f!Q^͍�Z�0WDb�?Ǧ*~�Uf��?Nh�浂(�%�;[60hPޱ�ܾ�@��@�E�N�'S����`�ъľs�)	�=]Йm6��ψ����E���F�����2�j=A�H��U@�BD���y���@c�>��ٸ�C~sL�0��ӊ��E�V�TK{��[$��(�K@�`���Cƺ�&�~�z�߷�?E�8�!�{���?
AF�$��4�'�%��\X�XRR���%mIӕ���R;i�_ht�U�T����~�{f�w��+��!\X��䂄�s_a�ȶ��fY��v�ƒ�	4�;}��-H��Jn�U/�z ��5K]��L�T��FyR��rs�3;5 i���$�mŒ'��I��TͅA�GU�Z�z�44�Z������P��ￄX"݊��#��q�������_��cޜ��	n%�S򼕳�w�%�g [Ȭ��嵟���'�� �7��e��y�%�}���Ï-�����4&�I�H���FϪ�������=��Rv����-�Tl*��S�ԩ��8�׷G��E�bː	�y���6W2�"׆���գ�jS���E,}�>��� � �6L��كna��TQF�����1�=pE]-�şF�3;���:�����RFެ�a��0?4��y��9i�F0������4l�|`���,�F<�xIZ���FU� ��L�����6�t�tS��ל���N�����@��*in���x5��v�E~��9�ASo����{[���>�B�I�l���@F����uB�EX�  ���:O���D'4,��E"ӿ�]�!�bJ� �������1�Ң�@7д؟| ����Nb�l���_fEX�I�3r�^1�-yH�Y%�k�-�UH���M[e֍�d�Yׅ���Δ�
@�?N1sR[Z�@?#����u��$.�D��S�}�
���ixs,�-m.q���I�uQ�ʊ�,�%�8���6�4򔬫��`�5j�B��ȧ�L��i�9��#���&�2�=J(H��Ik��Q�,h>�z[�	��k�$���Ң������B���X" *;X��|�o�q�ĜN&��X�G��"�>o����UNa_=15�� vBI/�tU2_YLD������ђ ����=�?�Z����f� A�gI��~�z�92i��5h;��O0\%�2E�%��U+gL� t�U\�ꉟOĔ�%6וuz�'�� 5>Ϧn|Қ>da��-��/�sQ�8nMX�:mG'���m�K	��J��W�(Jo}8���{PDf�����CO�O��_j܀&�`���+�2��������:��p�9�����}�qNN��I���[�&�[��e��r
�[�2i1��U6���do�4N��гhhv+\݅`�r�W10�O�4���"�_�P��A�v�X� \5Y��cb�4
��=����_`�?֦h1�����T;����3��0K�7!������G����H��R����������=dc��p��,��O���H�a%oZ���'�)��;;ʥ�����-
=��݃�@�]�Ϋy��:��V��ϦC�6ˠ�P�����7��?��u�:¿)��.��uB���Y�2���o1�}�$*[���wP��b��I�AJq����_J��R����鱻��T�qS���~ �&d�{�و���y����"�ǻ���N>0z?� ��� }��-���6Ѿ�s�D��b95�h	��<�A�F��$� �(�Rߑ����E �W�6����>/R^T��ɴ_P0��� ��'�`�j[�l!-z,m�˔���]�d�LCh�������6����Ӗ�82����j}�&�����?�˃肘�#��J���_	����:�����U����92�'���e��c������l<���_W*ޞ�W��	�\coȭ����l�R��ߝ��^���D�u�P�L�Z�D��&j@N�7ng��X�69���� ;0\ґ�~zC�M�_�Nf�e�=�8��16�g
�ύ��)�od�+"C���l�5L{���SN�@��H3fE?����f�I=yb0�5��'��\#�{��ϕB�_�i\��_��IL�G�`���}�cR���k,��ș�|:�l$$�_&rfא%ǫ_y��ݹT����jk �F-��**%��	X�
������Yd�$.�jBhVW�����^��,��v��ʰ�[Enf�[�z��@��~��o�P�k��a19J�ّ�f�`hM�tBO�K����sM���r�L{ �^���$-������]�=�݇�Ƥ)Q�9۸����6���c3�o�~6��J��ɕB�.�5;!���o�g��4��������){�<KX.'��6�����98}K�E���| ,�j��X�qQ�/bO�U;:�[�|X�L���Jrmh�XJ	f����$�6��>��J �o  ]p�~ns!*�}��T�>�8��v~�Oa]�e?���	s@�P[��&1G?,`Mq� G��(ɕ
�[ρl>�����Y��;'���|���� �"�6b~�Ak����˷��-�RK������J��2���V�{��C��v|�5���L2E�N��	J�|�á	=>���'����� ��cR�
l�1�& ���	��i����?�T8���֏ڢ�V��:�� ���cKkH�Wu�.::Y���W �8��E��w�〇"1>�l��g���jR��� R��*�<�lN����S��y<�g���(�7<�^�>�LX�ɕ��b#� �1��B�a����0�J��֗Ӝ��ҳ"�P��Ϯ�
(�*�']޹GgT��&���ẋ�Ϟ=�.}ے�h� zz�v��"��8E�aIyc�*��ݻȹ��+�!(������+B	(�8���7�í�ҕ!���f��K�P+��??��ɝ-4F�Z�پ�>�j��!t�B!El����=��q!������aٸA�Ya M����](���rr�[˛�\@����y�3�%�<;	�F�BBI�a�q�N�_�_fK��c0-k-c�S����|L9'Ǝ�����Wi�� �'�4OKU�Y�D�%ї��f��#��A�L�b�oν��M��}��tv���7�V��F��(�8�K\��fEs^�}�R��������a-�,F0�Cc��y��=�_*�;��˞-r��^�`�^z@_5�,.TlY����w<���]$��@�l���^#��.S�2#�^%X��ԅϨ�����
&�J���U�M%���� H硄�n���θ*C�:�`?9��Y.�ώ�����_vb�̤�"]�]C�܉�
VkG'C�S�6� ���4�(����qՁ\q,�%#���*A2͇��1*2҂�~:�q��~+�s����߆�O/nޫz��?#SE�3�
� �kg竴�x��~����9i._�Vٜ�c��U�J�7�YNԾ�}X'G�1�UM 1u�LOu_���<[=���a< ���i1�����4�
���29D�RVR�hD���˗�\!>��H�;!�yͻ��3�M�	|�$��~�סs cuh sjy�`��9i���A�`1������S��D����A�� *�9�Es�8f9��i�IiaG�ь��4`� �����9�3���ϸ�"�B�(�Mbt����sP�[�@�KK��%v�b�����ߘ&(�z���e����J���I?I1�;B��:y:ܪ��S�0�2XJ��o�p����IXw.�E
[���.��[����:��W7A�O��R���.#��0�m���D�zW#l:�u�8�xM�k\���4�VC_��( !������g�2_���"w�n��AAt�V�*�n���M����+��4���B1��7̪�mV��(�Vae�Z����3u2yw�=񙌊i��里f���O���f>K��#:ҝmT����ǃ�0W���H���!�mV��2l��s�/�E+`�^�0w?y�ɮ�\�o�J6n}���$�X���I�*4WT��V�{6��f~.��U.�����)O���~][�۷D��3{v,�xnsg\_��A���|��kO�>{Q�\�VQ34j�������gZ�WOB~:���8c��Z�!�7=%jo��O��w���dG�,U����YQ֜��
gv��6]l�t�Y���8�$�8�=���4��>i���`��o��d�԰"mf}Ka�R�h׫�xDc,`�N��,���$�8��Y�x�u9rC��ϻ"�F������,#<�柍�]-�U���#}��.=25S�!+������p2��\H��d�GK��H���.�^:4��[G98�3���QJ��W����Nߤ�a���j�0���|���c���|�˓odgy�N hPѭs�\Ob��6�1Yz�<����*��E��mH�e�<�jAΓ��l��531G��wc��N����;���_$�|��8sk��nX��^�@���a��ߪ��)������D,'�^v6F
��x�8z���*��󾳃��tD(3=Td��T�~�Y�av9�c[��%��+�@����ߑM��j*�����3jBh��H$����x�;v������^��}D�h�睮ݏ�Q.�l� ��!��!&�&���V �B����L+��U����Og�Ǐ�{4%�\u]4��A\���k�)�S%9�G��Z�dꈬ1��Ad�`�d	X�=�VEO���?�)��  �c���~5�xʮ���c�����$#������?�\o�Hέqn:2�]H�ڊ�t<"u�j3�����]�1l�HT׶�m�ز�o4q�ߚ���^ʷ!@�_�:?��^r�q����n�Xƫ�œ?Pt��:ś{z5��Q#�����"�!n��T�F�~����w7�(r�33��	,� ��9aӋ3-u��/��"�u%�A_��[�Y���B��zg�z>�!�wyIc�y;����;�B�IT�J^�3%Ư K�Q=�ߪa��f� �Z;!U����q8�ա�j:IA�.�Ҿ���;r(JmM������tk��2/aKL6�p�46(m�܆�yLz���U	���U�-�Z5!���[>s�ɖ~Q\�/����r��!Ƣ���qMg�7kʲ�t�D(_F?Dٍ}�׳�������L�6�L�b�x �m�0�`%P�!j�W�.�������VivFǌ� � �z�yA`�~S�	*m�o�ƪ�r~���/dB�<�DO念��ad��[µ��%�4�9�-���ҧ�
���xpM=��I�oL�P|��N);TTz���mj7�&���lA���\A��/%)mꪭXi��k�L�p)��J��e#�[v�X89&s���>��+���X��դ���	����hl��*l���j������g����];&ma��lQ����C�(�`jj:�	��ѥ�l��($"�b)��lq��˝�!��/bf�ԲX��r�l�ΡI=��r]h�lY�_U�+c��{?�L�NGp�i�	�}BL{�;a<�e�y�9��5�6:#��0��S26���Ε�)��fM���:�����NB:N-�E�sA�i̍h��ɲX���oj��I:�
z�)>����47�-]�%���jg�LE�3LW���� t�6L$\�Cr��E���Z�Y�x�#���#��h�䮅�H�,������ق�gOb�LX�ԡ`m�H��l��&q��
l���]U<��&e��	�/@�G�/����1��wXT��؏2�u� }�_K%d�k���p�
�y�=��_�/eL��g�jhzJ�HL�K�Oy�j�VN� �;���_���/�������8<�u{P��)�&����1%��C��8x�O�:��6�8�{�q6�H�w���Ҹx��n���v�e��㔛4�Vb]�� `I�I�%g�%����^������mҜ��oĞ�T�j �G���yNЌ�s��D�i:�پ�#@a�dCj����)SU�gɞ��k��D�Iƪ� �K�<S������5�b���b�c3��_G�IO�[M�h,qOiN���ֿ���F�U��T��M,���2r9�*獅�F����^��bd_�82F׍k���K�i���m�����L
"D)���;���OW2HL����{v���g�B��_�fO#��娗"yj�~7Œ�fw-�>;zT ���&��s�gq�
�B/7�oY�K����K�F	G�K��̈��ӚHh��`��L�).�"������J���y�k�/5����qt�F��C�T#OV���MnI���.�_��>��㎣�8��Lֿ	)u�����>�	S�H��
6���v(XbB�Q�sϕ�c��C�'�9 Kt kKk�Y��vZ;���CB 1�l��\"6MFޣ��aW�+���J=ef���(Ҷ/�1{�o�Y�L��w��vğ{�b��Lux��m���|7I-vs��T�	��'����%4����j6* +8牅�
�W ��+g�����v�:�.:JZ%�~�Jp�� ��Q}"8C�u��H��|�=�/BL������s�Sc��X�r� ���8<y�]�/��:^DP�"�P4Y�I�}$*l�Hq���
;WX��l���RtT0��u�AW�Z{��l�eI������3�#)��}��H��Ϣ`L��� ��Hn	�s�}w����
�fn3���&��|�O���!蝺(<��8��FĞ�~a��1��RG��
~������Lx���ۉ����S/"��|��T빢����҈-�_+^82ȇ�-sg֊��fb9.�|	t�Mk
�I�M+a�Z�q������X'pN ���N���V�z.ڏb���%h�nƜ��(VX�� +Rl{��(.|�:gƪ��[�Qm5�M��vs?����f�U�,��Y5�%#�d�_�_��ܞ��.7�mq�w^�� ���ȹ�1�2����p'���4=J`�������ʼ���LTx��T#���@u�P�x�F��JF٠'�Q�f8�ϧ�q�/�a�����Ӥ�a
���y�,M%��`�%eD3�J%j�]���ѣO�(���Ж���?f�!�H!�J�Ut�X�*J�2�Xd.�H2*�@MHW������Z��҉+"���������H�WM�L��ǫ_C�]�}�q���k�X�U��n?��7���`:��|^��P�CqF[<�[�B�Å>��;�j���f��"�BF�n������,釨���{��Suͱў��'4��.�N��}.Ke��^xr�s�I�<:6MK^��0&E}����Q��A�S�cr�b�dA6i�AR�ü~ ~
��'i.��:��n�Y@�흏iO\�B��?�x5�JI�_��E�mgh-�4'XygM�xOGt�V�S�������v��;垶a�'��ܩϡ��A)~H�ν��K�bN$48�(頟賒qVب�	
�����Sh�`,���!&tŷ�c�JY�4XZ=ǖ�"o��Qb�>�i�R��vx�i:�w��<J�! ��¤�2��c�r*O�A�06�6�lv��pՑ#C�WE}�Z �'��Ai��U	K���=1���f��>w�M?����k@���l��B|0���uc"n'쒄��g��m4�.�,���f~D��u�MiԾ���w�i8�-�@-R����2�[NF)���>m2��]{G��<U�m�i+a�-��ȯǮ��=y�Â�����vц��S�n挋8�'U��y�C� ښ�%�0��Zۨ�mn��xJ�4��.����� =�)��^�0�5��@ �����iH�]�=�]e ����I���0�S�����.�0~�X�b{ߩ<-��$6Am�0m@��px.�s�Ж�o�F\OS�#9d�H�De��z
d�"x�8횓�S�|D�YOT�1ͥgð��J�{�a��?n�%�����A�Pr�0=D��3��\KN����T�?�L挀^���=�I�R��l��\j�h�S�GF���Z��e�ݟ.j$;ޞ���a�'�'�3X�&>a
]D$=z|;����;G��µ�Mc�@d^��]��l�G �/p�"��f�cE�3���Ԙ��;�l�Q�ll����܁Fئwf�����TmmaFd/`Wٶޮ�\Z7��!v��	��\4#���f�U
���x�*_Z4^��R�31Ԝ��+0�����{�
}p+lTA�&���(��+RtS�9�2�tZ����d�k�X).�m@�%���kʕ���iH�?p�� �����K�x6�����_�l2V��=餢-�=���{�0P��U���>pX���!���Xݗ��0aZ}�m;�*Y1�'m ����r�5�$����*�۝i}� ���fF0��W5����lU(5=Ԑn�i%� N���/�7��[�Qr��d�v�﹗�,�-�����eu��z�%���4����Xu*�N�����7ٔ22���]K3c���W���\���r_��UV���E@��PU�a-n��9�.�����*F5d��R\���)1Y~xَ}=pL���جlkh9&f�o��ǎ���ĪCk�n���X;�19>6;�9���rop��b�	��戏6�6J�0���SZL	5���c�4�#�DuBQP���޽����	��0B�9s�~`7��̳�P�M 3*_>����~�j�L��`�&�֑/P	\u-�0����!uq�N@��������MN6yG	O^��ګ��""Wg}�< �oy���s�(�����柵A@-����`	wy{���oZ�Ŵ����6C�R�m}�C�LW�)��g���rh�l��[Z��>�C�'�뻱ȷ�"II0D����h����� �]����|'E���W�9�Q������ٍu��d��S9�Bە���0���K��W��9x?��k��Ls.���$�����t�I�zgu��壔��z�?�������Т�s��̩�V(n|#�+)�0�e�7`k�\�k3sv(8kB��-�W��oM�	�=d�&��է��bG^��U2�rG�U!��?q4wC���d*gF�+��i�=H�����9�d����)��-g���o؜���Iگ���jLPw#2,�ԩ���¬`����K�7�3O��l	vQ>�Ji��~�MZ/�3�i'+�i�9�7�D'�Iײ&����Ö!p�8���s]���\�)�+xI�(iZ�(�z^%Ad�D��R��pB]�;>v�6�������o��j,,Ô�N,?��G��b�+���`�f�H������a�e�a��4��e����M�_���Ub6������ ��F�Ƕ��=�*��پdm��,������o��su�a;�]��2���:��\p�A�iɛ�1NM�����f�&����6�����EqD�o.M���úN���������<�����{>&,`u�y�&��+�3O����� +�\����q����xe��Xu�S����0��vym�ؠ e��/����fi����j��f��7�X}�I�`�<336�L�Y�Vq[ E^{�r����)pZ!#�\���`}J��_��	ãw d{',L���ôP����B��}?�7�X�w�jf�JǄb���k�Q�@�������[W<��](È�&�OoR�>��?\�Q���|�)�!- S,h�0��&_���5d ּ6�[Q�-G�1z[5֌
�p�8��1v(���t�
��rT�&o�$h��3�e�\6a϶A���m��T���)|D��	�;<��0�!3Ƿ�t������F����\�Z�X�dK����U~o@w��Ћ̵����O;�AO�ıö||v�H��->�����@w=�#ݿ�PD�a�i���L+f�b����	�v�fΝ���+�Mb"t�q���gf�j���c8���0�A�O<�9�i��G�G������� @K8X%�
S�Eϕ�C�>~��ԅ>�8�i+j�P�5��DU?.�� �$	C���<���5h5o�u�%e�^Qr2�<߉�����⢴_�w��������l���]c���(�-��v���#���}��>�rW�oi��
�S�O@\,�>޹گ��V�v^�]G�4��U�5�ʖ��F(i0��=�踶�ui�����3|�ls���^�ܹ��f<��ߕ�D�ϫ�~�Z-
J����4N�w�їxc\M�i�$�wl��GZ��8ˌެĚ���|*�2�ݗ�f��7ǜa��k9e�s��#.E�kG6���Hťp~{eYVE���wX�����o�r����!�\���)��3���s�M��r$�u�Dޮ���v3x�����c�z	���}y܎��r8ud��l�z�#8�M� d�ʷ���R�A䲙���$����5��uoX�sL�,�@^|$T�es�7� ��Y9@��7G�WZq��͊��I�y@��a�O��/w�O��<�z�'���M������~:k�]�C����'M;�)Nfb��pc��O�
�[�'��g9�2�2L�u��5&O��X�]i ؁�]"6v�2��%�g����3�Gڏ�X>�Z[�Ĺ՜�8�����R�O��o6�g��h�����5�<���ߚ\�i~��§�KT}
E����-W�x3�g�;���%=��Z�>eG����P�[��.j���v$���^���bˬg-ڐT)�:HI�ʦ<h�N��G}t���J̞̚�X@D�&���Q�7��4�ł:u��8��Iy.�C��T鋴�Q�I�g�oFO�}ߣ�j)���2;?�K�*lv�ԏ��@��;v+�<�������¸R�ut�w0��(o�~�vu?�S)�����[я|+j,���/b��nv{iǢ��ݼm��-A�?�_�Jx�SAE�܌�~ZN�!�_��ݔ��q.��	�uD�܃f�!=��Z��84����]?��9^{��Br1Q[���ù�$	忚Bh�OZ﹘���2��P5��`L�@�@��NO)r�������}�|��F���X�~������/3�4V��+:5��e(���6=��f��E��p�e>�ՓDգ�p�,*ͯ�j�rW���xUa�G /�WJA_��� /��]��C�^xj�8�?� �`O"���p ��tkvv����
�y�#r�8�"D�ڢ�#D�%< J�%��%f�]W\x�E�)�T���q.f�8�b�G;֕�Z�P����'ޱ%i����v>�I�˕sTys^�Z��m�x��5�/��A�;��z�d��Z��5�Ŏ6x��=n����������F�_��S5���C(��+&n�as�n�c�Q��n���d��7���Ī�iiV�5Y̬ ��n3�g?:�c��E�\� ��vo7��($᥮]�wݷ����Ĥ�A��8Y�aj��]o_��2p�y���mH�!֡qytG�]�6JOm���B>�G��y���%q±�n|g����E1�I���5�\4�	V1,-�s��qfpn��l1�B n'~�\�@�����L�-�� -,ްd7�XZ�#�X| g)���f��j���V�9{�	�n��$&jC���Z�-�o'[�x�g6�"�7J�5��Rn���H6�5*p���!%�8�>5n�K⯈$�� N`��wLZ�3]=)�D��C��R�;�r-1#�(>~O.8�~��\��e����h��&��Z��+Ԝ�*����5 kpK����4����a���-�.�L����?�F^�d�� ^����![�w���B,�2�6ՊfG�V	�zф�K=^�:�~n�_�������g��x�+��4�]����K����-�����x#��	�M�:W~���c;�XP^#��.PLx�09�i���pj�o�Ƿ��h$��h�f�B���AX�lӞ�f�ɏ���a9E\��`M�>oM+!��R�A1��@�.H�f=O$v��X����H�
��<�q�������Z>�	q��z0C3��)L�pX�ndA��3�@��i�=�oV��}��X*dB�[�`���IDۺ��c�����ϓj2wQ���
��O|S�0�����?L�!K�o�������m�P�R�_
zt�h+�h^����EtՕb�R��]b>�~^�PeG61>��9�5��9X<�����`�y/0��*a��m܇��� *��%rI�Sȷ�P	I2Z��a�1VQ�W�5�%���*��0c�^$X�Vʕg"w�<{�P�9�:�,x@Go⚕���<}���~f�����7�R6�H��>�� ���$;e��OLz֩.X�"�t����\���"?�C�Su�uQ���� ��R��2z��-�Î{	�^�Q���N��q�e�8���?i݂���a��gʭ���w1�B�������F��@$��g��3��s�rΟ79X����ת����{�}4��6�Yt`���D~J�Y?R�˗�l�7FH� �$�)�q���2�t�Ik>i�uI�8�#��%��p����iWڶ�l�X��F�B�J�?�M[~��Jkʩڗ*?uҝlf��zT�؅Q�:�����.��X�SI��&E���܀?꟯ ��b���7#��/��Dcx�G�����<��X���v�`������4�w�1ӿ5�9tk~LS	�8�O�k���A`UaļL(��<�q��-X�̈́��V�&N�K�����w��|^�L�?�Sf�UYyH�V~5lY����_lM���T:lʊ�-�"�����Z��e�Z��.uO��7b<�r�	�`�>�7�QK�i��!��Z]##QB��70[�K�CP}��\tU=+`%o�;G�h�����m���2gT!DP[���$"岧���ujhT�s,xI���+�G�� �LqS,B�ŏ|�eܑ�
#�4�ng�t����ێ*���&����*�uj�;%�m|!�t�#n�uS���j�����*��=c�N�8�h(�>�0|,�5��&}��x?��ܤ�S�0O��%�����k���X0��E�D�9���#o+����5����6�W��5�E�ɶ@V*.C�fvZP�A�_Z�E1��U�z���+_fb�����<��[9�>�,����C�'��������AP�=�B��A�K養46�~ǐ&:���c[E�w��NTդs���J-�?�uh���s�	ǒ'D3nq��K4�����I�ԛ��	�UKB�rB��zE��98ƀeM�yn�g�[�{B�g�;���a�22f�3����3���r�}��#���2�xC[3��C��T�QF�v��Y���v�V�lE����i�>1kd��g#lfh�N�!Pg/�:<�㺳��JȵX{��ihf!_�ۺYk8��E��P���eߨSl�R�6uc���_=�C�+�5X�������ǐQ���5�����X\�k֬��/�u��U\�aV�	U>��Pj@�����~;�p��6]��_�8��=m���',H~�NC����R�6��/����ی i�i�>� ��v ���
�b����xӧ0T':�¨ܧ%)�^���}��Wc4�$���D�#gw�H&S����h}k�x�$��8�x��t;H3h��&o�!^��<���W�b���=M�>��jl�@��1_��7��?�&E��FW�B�^ק�0Kp�U�%q�Z���i&�!���m��.$��F�aӫ��6)!2��%V�[�eH-RD�=#��<�wVl*���)%'=�;�$��R��Kƍ1R5���o�9��a��� ��l��F���̱�g�b�|��ͪ�+;;a6�D߿�r*&��4�u���f�(�y͇�]��{w��p��*n�E�-��Ө�1M��];/��i��վ����6�x�(����X
��r	�?Sd ���Jl��n]A_a�����v9��UP�N��#�|d}H���_��ή����ց�r�j*��˗=P�.-ÜN��ld���l��������k�4����:��#t��h��G�:Ek�cC��J�~f�_g�1 �^�q�����I�ګ�c#�g�9Z�RA�������t�C��_��5��AF��WbF��j�B������,}*�'dZ�����Ɖ���h��-�5�ZvuJ�S �XuH�
\���#�n��N��j%)��C���Z"ݢ���D�,Eܙ�?��R��?����^1��;$AZ@[��o�{���	�?�:mGIb��4Ww�c�c_��-��N�^�xb��[Rl��bs��8��(}0)���k�p�k��q����0}: <��?HKcJZ$�л� �G��d�!��f/>� �2ҙ7m"��x5��:��+�;<ʪ4L�8DÍS�C?�BHDak�O�%�@V� ��b�1��N� �������9���r��b"�ɯ�6J��r��R%�.���i�deg.y��R�sg���+8����K��ێùJA�f�O��)9������u���U�Y�Ɖ��%8!�1 ��?�[ ��� ����e1'.�*`��K��qB��+��j�:��aS��lm��fۡ~�Qr���K�P5_��X�_:�xJR���~������R��R�8044��,
Ke5�m����y�d���\7��/��!�dh�%
�0:؟���pV�Ы����i�����)ϴ�@��z��;�Y:�KP��.�8�+��IփS
�(���v�>���4Y�A�3:?��w9T�&��'��%�����㓒,��cETj�yp2��{����хi�ICg�#X�~/\��`�3��v����O�A�L
�����|�Ga�K� ���屼���1��C�Dj�Ěó�N4��Zc��	�>���:��oCn-uEÊeg�.o-ލw��W@S�{�n ��H���D�:��ƧVѷR$'h�K�8�l~����m�3���:�?�4���l��G���.���:�����@A2>���;��L��y��K5a�a���Ə��̣�feK������f�- ,��Z<M�k��/���.�b��[�,�K�"�}�Ыe}��@�����y|�Gm�s׬��4�6
ħTX����#9�3�L���Y�)@�p��,H=!6� ����G�L�Ui^{)�iqP��������S*��p0Z���ADLT����;]AJΌ#��y��Tj�}��L�ռ�^2 QjqY��}fB���#w����q��]@g�*��h��2	�0�L�'JkK�������2�暎��ǭ�E7do�'�*H�s�����{�I��z���`�J!z/X���#q�Z\D�W�6���S��b��Ē����`b���/�KBa�Z��\�%X��Pɼ�,���h�c�(�q����/�E�-xX�T�7WUđ[�5����-|�Q}������0(v����+��]��3C�>��Q%MJ���WP}E�����V�^jiF�䓘����z��O#a�t}R{ش�ϐl�ZW7��/_��q����C9�R
�B)�G&88�/c������7'FZ_p��:cң�����(T�,j�?j�My:�wh�#6�8�� q�qG��i��;&���
��V'���Vw���(���i8A�З�h8�_n���*�r� ?N*�J�u>�o'n
��"Ըwc����	P��KNهl�Z���+�c8:�6��ǥ��n	�E%��A
.�b���|�t ��[v-���;/�W��7A�,	��Q�H	�ZX>U��٢��[�?�~V���m���"}�(�IF��H��A��ao����s����i�����*�L�+5ǯф� r�Qm@��* ~��@P�Z���ߓ��{���3� �s���¨��N�:�fb����7+��H0���r1�~���0)�o`5��m
�+�6�g~~�x����Nۖ���o�C1��*�".�q�jg#V��v�v.B� W����e��)t�t�:R`Ι� �]vZ�X��d�%Oo��wVI{)��W�S!�^�R?��Ƞȧ���8��I�T�;_��g��-��0"������44sɿP�aG\�Gq]�32gϩ��I�˾r̰��Fl����8�c�&s�7?F��lm��x鞍��tX�9�97�ZLN��-u���#H���{��G�l����ޟ�˘T���2ł��� ����b;*��L:�g������Q�)P*�]��Ycw5C2"7���,y8�g�6����j��蛧�a	ف�_k�B_q	���ˢN�@�B��/�	����fUnЁ0����������
c���o����+�f�y�Op��k��
�E%$��@t�}S��+�Bm��q�ntX$�״(��4������wA�E�~/d� ���i$�QX�&ߍ��8GP �écN��*�{�1j`G-��|��>�pC���SL���C
��J?�|Af�s7�o��2�>;���) $U��pb�tJ�uT���6H(|x�_��aӤ�Ra����{�oYBC���d+b��������]�@:���f	�^�Q*7�/� ��. �a䲄�$b�k��헩�؈�6#�3���l%2E��d�M�$���P���0��}9Q{�V"�U
&�������� ���l�]��-�qE²��#$��
;�	$!�7x��M����ZQC{M�CH{�w�Ql2����2ǐf�\HJͶ���@����M�fV8�@����ĩ{K^v�4����s��M(.��i���>�W���}u�|P�׻��}H��8�{{2���պ�fp�do7u݋�����C�1�w�f6�y�E��Gyj�d5��P�����U|�\&Z��'���Q���2��(9�U�������s������W�&��,��p�9��՜�
KF1D#�-�]�țu* �ao;_�~D�ꎥ-C���$�M��_0K�>�P��И��΃o�������������51j���u#X�Ut��,�Š|s�p�PS�(�o�-�U��¼�R��.W�A��f$���n}c���R�t�̙݆���
�m+^s��FݝdH7�?����բV wt�3�J���tjw��X�'�| Y�g$���D:�S��3�2?�R<[LZ�@	{0��[K��4�;�db��%T���A]��H8۠��D�o��F�4t�/Ǎ��9��-9q@Yd�n�'0�M��~x]?�1�5�x5�Mn(�g9A\v�N�N2��\�@��D�W�j"���!O��CJZ)|����_;�o��wD^�7�ưUC���U���	F����hA��>w9E{�y޵%�0���m�Q	�uް��&$}�D�=v&A	h�(Lɵ�-��0Dڽ������F�%'~����s%�{��(M�?�Q��#~<���,�^��ӭ��گe�io���ƣ���a��
�k�U		��݉l�U=&�ǥ��J-��l@!�n�{LS�N	�#��H~�m��H�_,}��!&���I�f�#�s!I�c@-|O%z�����V�R]�B�.0�V4v9��HY�$|�6�>�jW'�*��$l������y[�5P������&w�Z�'�}ĵɀM���wq!�wq��i~X"��,RAO]���&|�0���)��<y�"�a=z)2���J�*<h�̈́D�i��o�M����p��@�O�� ݇��,r�wwYJ����Q��Yg,�Ku�X^��)h���t񹴢�)���{0�	۔-[���s�(�h	eyp���OB�M><�����˪z�~y��#ic*�a�nL�|��_�uY�����6�u#iSB��(׎z����"�tD�h�`"֯���Z� R���x2m=p��@��z6H|���ۡq�j<s�F��}�������F<�����n���|3q����.nuU����ᠹx�c�����8�@+�~�T{�^o������CO�0:��wJf��IYv�|��"��) �h�I�LwHO��.#kŐҝ�Ti9������`UٱP�>�!E���>��^�fl��o��Y`��u%3!l�[�q�������5�6�%��H*IO����b跎b���S�+��(��f�l|��v��ݞs�V ���Q1 �&��R�j=��T��e_X�˺C ל-x��\�ɍlF�rn����
Ƭ��P�bͤm�P/5�DD�q�ϛC�����<!w����A���.j���S�w��B�]����W(x$V�'�Á1Ŀ�
�P�9���(o���t�6�n=�&��C4&�Mͧ�����J�8��U��y���NB �@y�C4w�!��S�� 3:X��4)+�]�R�a6�a��KU6��B:y��	{5
�~ÃY����h>�7]t�;��`��X��Wi<�ۇOܶϯˀ��}NVU��W;���Bv���RaV#rfI�P�ٍ
`�ZZ��E�m#y=y�J	�]�,�JZ���(O}��]��t!/Yj<+7�&�2q�r^(�m��B�[X��� �:V�'�� ��+�)����5��(+����YF��x����M�����;�"���w�G0�ǠP���T�.�C�'ۆ�am�s%�>����FPip3���<��|��)�!�^�OC�{k�G,{Y83���CьC=d�\�E���Z�����E,���Rm�9�겵;sɟ/���������LU�j�5@@��RD����쥨wLJH4[�柘��R���Z�i�L�NE�P��l��Ԑ�ࡣ㇧;T�@�7|�,J'Ҁ ��G}}��7�^D0�/τ�h��03�� ]���SV=�)���g�$xA�͓G.������b�NS��54b�Wa�/���E�s�e��f\8
hY5O�̬N#�_T7��I|o�k�1,rT	�Z񁄎:v�c%��\i.H&W�\�;;���?w̳T{$��ZPT���Z���<6m�Z	�:����z	 >%���e��`JGŞM���?&r�m�f́�C�O7����P��0�$ǜ�l��b	���qH��&�*r�j�����m��.Sv���PA���@�R�d2�3�D:ǹ���C�G� X��'X,�u�hb�e��i�'��K�aީ+eS�4���X�gkbh�6cQ�rr����7�@�'�:�1B�؜�`���=G1�j@�t���A�54o��NH����Q#i�g�2�&K���g��bO��*�-�ܪe��M�%l`�>�� ����I'�96�d?���V�0�`�G�|O��u=+�%- ����,��I��3x6P�=�ΨӍce�=�Hl]�9��wѓwB�:ꦔ���[���@�%_��
����?3��8)�;��?`w���?7����ߘϻ'qQ>!���v%fV�uֻ����i�߇����x�Y)��Y����Vo�Y�>��w���,-�@�����7z�] ��Gi�J��e�iG�.��sî�6�߲�m��wr�2��΍���'H�&W���J.ܓA�[Ĕ��XYɔq����!f��B?as����A��\�+���	`*\�+����`K6�kR���O!�k`g��ÇBZWk���wg�`��eK�K,�J�q�0� ����;���8C�,�
���h�����'?�i�����U��ڶ�x�
u�W���5���1{`Ѣ�is�%-斸j|��<]�?r�Y�ŭ�~J�+(y��0���p^�Q��6MI�m�N<R��k�Ǘ�w���]�=�(���x���ߺ���`��TJ����jT�]W���Q��r�U�����O(n����o�IBQ���y7#�:RΣS�N����|��W$0��9�8�c\�mu:A�v��i�8���r�e
b:�>W�� vDG��l�RF���]
Ԇa��!�~�;ۀ�ÊZ˝�,?�g�Ȇ��/��/ǦH0�'szB�k�^�oN)�:�E�˔�`F�Kk�\]ej�W�o镟�^ �YO�8�����2�{��uE^��I3(l��}T��(d�QX�_��X���~���-�
�>C���g�`�:d1:N���-�&1�_h|��]n)�D4�J[$3�4��7���j�IO��F���������Ө����RD_	��nz��2�r`8���}D�R.��C�(�����YG���}�27�Şw�KA����t���߹�h��{�0F��"���9��+�%�#,SղyqѤn�0�k���n-�cvy���Y�O���̵r���|ZX�F;�]aLZ�PmZ� �x'�qn�B5f^ �ٹr��Nd�/K@L8I�R�s:�IoB]��=1,㵘q��׺Hw�j ����Z@�#��q�b����/<�q8�u-���ʍW��=9q�a�(�̗U����%d�v]X�l1����.r�w��L�nÂ�G+/��S��_�\p���VN���!А�N�q�NI��ȍ*Ө8s �hF�x��=��Ǻ�ze(�DB�N
�� tdI��_��O##O�};�^�I�p�oW>�3����/�54~ �,@=!2��{k����	�)�p�G?�3�!K�֟8K�Ǉ�	��L�h\+S��[z&`+/��"Ԣ��_O[:"j���̉uD�H�tD�p��4�яLap-��%pK�{Ⲃ��4q�U|�0NV�iZ
S�p��|| R�H�h^�4퓜�i��M���\C���r�3�l��cĂ����'�C�n���?�@��<J��j�&�ʹI�S����k-L>V�V��1G+��t'I��D�4���9B-M�P{�Q{�_�=�1��h�"���3ܛ�O��d��P�Y��+W�هà��c�y�ي� ��=�Gh�.��<����_Hcq�mZ[C��]g �/��v�F��4{���6O�a�;����+�"~$�#�8j�6�1=�Ů�?�>`����n8�g�Co^�`ĝ�|�_zS�d�I+	.D鮘�1[<���Ub%͈�$��&8�!�K��䳋0�� M�g��T�#�������దt{�iV(���>b�h� ��2O�s��Tu���p�Cb@��ҹ鎋a\�ޏ�c=dGK��P��֩�$վe�u�jΔ5P)���b�\��;����c�(o��瓪�b"#y*l1�[��ߞ��jMʹC�n���|#,T4W"tL0ѷ�{s N�����5^��5LUW�tR��b��	E���K�а��Gg�㤒<�.J|�g����\ͼ��������q��{�lv8�(�\9v�NO��,q)��!�w��b�ԇ+NY����}Og,��L��*�}@�����W��!����o���2� H�ؙ-�Em�TDdve�&�E��Hʳ�����¥���~�����rL��X.T�8y��:O�{-�#.�3�;AZ���\z-4���kފ�OV�V��*����T#z�}ڜ��MW�g�V(^��Tb�*f�<3�������}�<����S��c����sK ;��
g��py�)�������D��R"b~w�7M�-d�"p0������o=�T���^b��w'I�s];'���t�m���J4����ӽ��.�/��_�7��o#x��3JS~�,ن��71���dx�a�Z�����p� ੖��h�,׌w�*�(�N���a%�/�0}U;q�s�_����gi���'���-D?�����^���8R�_W?���p6=r�Y�wi=7��rs!��m���FS
��|�\zZ���	��cU诂�K
�E�d���������o/�B��2/D}4C}���_�˷�sHʆw6SԚSp:�?fl7t�S���W򈒑"<?�뎕��3��JV���q��Y��RV���>� �����l���|5��T�ؠ���;WnZ��JˮX�b�0�ܷ��P��=zr?!��i����0�R:��{�! 1��H�����3�V�l�����N2��n���p5l@p��dX�~�	B�������s��?MI�@g0�H�s8�B��G%�,;�I����)U�r����} Q��7���H2>S]F9�ɽ/zr��R��yd2��`��	�]�Ҧwk����"k�ʧ�s;z�D?��݊S�l(L�O�vW2��j_T}�� $��W(�Z�V���vӮd5��XI��={�:�7���� \��O��i�3��Q0J�qKa�LJfF����+Β���Y���?�&�1|��B���\-�٢^�HI�(`l����dk�2@m���J�I��Kє����r�KNn.t/H��n��n��-P�͕��v�M���~GO$ưp)*���j��Q!�h��6j�q���z�,�|�W>Ԓ��w�W���QB=�~���5S��3@̴'sO|Ƿ�`��l��/�Q�L�$m� BS����n��Og���$�L��&��[&Ճ�vO���
:��_�Y�}�.5j�/f�<��Q5�(C���Z�~�Q�ƚ��@� 1�	����ޤ��$�I��u�+�6H8?}�r�z�n9�]���E��j�D��o Ny������!"�)���u:�QԂ8˛�(Bj�J��d�R�^B��H��o�/�9(����/+OX���9�X3���Y���Ύ��`�4����7�³&CMu˳ ;����d��w�#��0��ƣf��"�S���ЛM��S�K7���E'�
eP������jJQzP�+~��j��>}�P�\P��e�ۣ��n�l8z�@*���Z��v�T��Ԣ�y�����f�O�-,�@�JW@�9�!��ޕ��b��Y��ӑ���Ι�2 ��AA�s?>�q4�II�6���?X0�T��rhs���O�s@�����0tm��}-��t><ȕ^�Q�ȉ*�x�+OS���gOb0H�u�Y�T��D�F�,%����	���.�(�>�����rn��|.)���q3�J��#�q�
{,�co~d��$ٯ|"��8�`�[�o���rzw�/��`#珖D��YH�l�4�w
\�v/YWy�^��݄�XPn��Q����}��Pq���O(�~�0<�;U;{t�B��wϙ�Lk�YY�b9�f��*|)�8�_3{�͑��$ס��[��S�L1}��Ą�,���K�BЌB��W�(�桫2I��8;�uܬC�yZ3��^=xZ�>�~x�h�y�u\E��[��7�N���r�R:�֘��0�K�Q�x	�d��coJ6d���d>a�ye��7h_ q>�,�k7���<Vz�mz��;�eT�%��h\ަ�Ҽ�lŊ_ԃC��N����E��Pw�ՃT�W~�)9�B��sg� ���K�F��-4|KȚ%�����͏��v�d1E��)�xi�rr��p4|�äs���G�i8�-:{��ey���1O/Dh��L�Ѩ}n�~�|�9�$B�	y�� �����f�H]��-1��C���.�A{w�6Cg���{��F��[P�?w����&�U;�"��:0�@��a�ś���<�[�����_�K����\b)��	�OU3,h��Q���?��432����s�p����e��;$xF͇t�s�ae:"o?�2�����eLC�p-|�g��B�`�`Ҋ���Lg����b�
L�{=;�!��j��dr�dz��E��C&�$B-�@CT�����
���3��X��S��BVaN�敔6�	�;���TU��Mq�1�%}� �x���6E;�۰�J-�ԀYe����$�FG=S+s�V{�򲉸�9�'d�J�.E2��KW���T�n��g�|�8�M9��7�ʭ��������[wC��Qn�ҫS	܁�Z����oA/�8��\[�N��mYr���������B�}��x�����0ћg[�Hz�.��:��Y��0GO�D�h\��9�P��N���?$�%��w��x��@d��z��~Fc�C���i�FE_
Yړ&7w�
Wd���m��6���1w�N���<��k@��aa:�(�9���ʹ�ދ�J4[j?��\��<������l!F�򵗂ӽlk��������^�3an;��l��D$en�eG�В�ht�{��N��zc�T��sU��1�a>���PO; �M%�؈�o6��u� �M7��v�y��,'��y�.� T�:E����!�?�e�qv�\����ih't�����r��	�@D3��p7J9Áe��Tz!R�;g���ËZ!�ʚY��M���7Hb��ލ�* ��$zR1R��32�S@6E�۾G��~Z��_E0a܂��"��y��t��ô��Y��jB+���A��J|����7�2GM�t���^�����<׼ɖ�^t����������]J�|�fly��ѵg3�,��
!:�݇�a�����F��l����'요a��ZD͔��~�aU��s/�`G��q[cF���k��O���G�V�N��.��I021F�;���&M����e�Gfz�1s���F�.����/���p�Jo^�
�U�~�����2=%���wB�f����>[�\����ۯV3�#
��N0�ɩZ�O;��F�TY;����;�h@�uw�H��?��*�D��܆�S�9!>�ܝ9�"�p(t�����U{�G.�ܫ��ik��O|c����6�3����+���V����k|��N}~��z�ٲoς�6���<�kf�$#8	ȯ��+�w��12IKy&�F����,�?-�e)����aH�kI��5'�Oa��,������$MS��ggk�
K���_׹
ip�PN����BJ��1|f@O�Ft���
�A�:�{q��֕U��pd~��@	ex����c�@�2�
��Kly���CSa��&�3���f^?:��a�_�5�q��ҷ��#(�����<+�2�}�j ��.?�&����g�e��������)ȃ���9���7l�m��]t�g���]�o�{4OV ��"�B�>��ȱ�u� �I��5��S2g=����D�s�&;��%\`�VJ�R#� L�6����p
A�'2��k[��g����̹H�b���)PoQp�J�Z��_�^�AWY(ޔ�z8���
��N� _7���n\����.��_h6.�coB�'0co��n��Y�O�״�+�����|2�*���ya�{H��	k�*�h�ō"�$.h�+co��@���ћP�I�n�׫��+
:m/P�tF|�A1���&ku!C�LҀ��|1��f�,]xl�Z�C�qpE�3�]����x�3G-?����tJ��M�G/�7�6[�g}�@��d
����D/�B�]r�c)�t�P��8��D����+ĥ�k'��<҅�|ص5��?�!�W�5�V��,E�X�h��\�Z����!6v- ��#ћz�b��L#���!�^B�^�#\��؇Jв�Y�u�O =Vb%Ⱦ�_]LMî����_���BxW������=�*��jZ�%v<�>s:u�Q�rOھ�6��ud���z�Z]ι@Q�Y�z5mP������B�*R]%J��l �Q�V:)����dt�z�E���6��g�Zkv��d�X�XG��*ԁ�Vϝ�mK�F0U[�f���	J��!��;K��3���-�x]7�93�_�$O�k�.RSh�H]�=�S�	
/���M~�]>���Db��G����t��$��[.'�s��V��\`�qF���n�YQm�iv5� ~:�0qrP0����KaEӸn��v�%]:�:lh����� �CN� p�v�%[%q�oy�i���u���4%&�0�9�d���w�˓,�����	@2�t���X�C�%4��^�Z���f]�)v3F�$G���<g��
Ĥ6!⡥���ny]gb]Ǌ�:,�+`�j�O��g��@�]���A��r2u�N�������5d- �GIK��Y���ȝ~$&�'��A�e��5��B��G�0�ape�*���
K��*m������rYٷ�K�f� X�Ch��V�q��]��h�bQ��[Ř��/����8I���3vuN�t��F��Jⴃ�rĚ���|{ƛF�1��1Kox�U�yN�d^C�:?�["���.&�r*ye�3c�ህK����Q�P HY�Up�n���ϭ1�������γV���6��չ8�FժK)~�If���FАƲ��b���3nR���
�Τ�҉	(�^�K��U��Q��\Fd	���G;D+3���E8(q��q���mlT�*EO�z W���m��H�Ʒ�+��kl���G�e=�ˆ*=FYb{H$�!�ܹLһ��[;ѿ���4r��MC���Yr�
��TO=���U���,��L�4زr�G��uB�`����M{̧�Ј��|��?��gZ�َO�V����S�U�P�����!�8�PNju���V[?��O�FD�X(�ĭ��aJ �zO�_��Ol��"�������Y����vg��.<���v<4͒:��n�`��� D%�󺘎�Do�e�f�aaѨ�"��a�Q��ؼ�g̩k�ܸ�ȹs�z=Q-�����|?�z�o���x�KCZw�j95�)�e�j����*DD��0Yn�{*�T�.qNv�r��;�e��M#�����a|� �c�\4L��W����"3�(N;d77�̍3^E���T�l$i���ĨE�m;��>�����=�*XO��� '��MQ�A��`�+�c�-=�D���m#D��.�!u��x�;>�[{E���]R*�'B"����%t�c|a%��M�K�����CԄ����~޾u#z+���e�k�N=[˸ @�:�6gr<�YR��1��Ao3 3"��Q'3(c��zL�s��z43��t�(EݝȦT)_E���;6��C`9Ϯ�����ZX�����ƹp���FAtJJW
~��]��#��,2@H�i����o��G�T�G��=�2��獷�^��0��{{^�L[�����؂��^ Gp��٧q�����x ��A�^5ɋp>����t����F.�a�]<�u�]��B�NK�v���$=�Q�セm���;�r>+�3�ʋض
|�p��^��,��G���컾�4-����:��Ծtm����ڈ��s��&+.e#���<=�*k5��6��u�NT�WD�
=}qx�q�-��EϘ2�ne�WB�:�d�q��t�E@�2f̲ �a�Ȟ	`��тz����W��f���'g�|rw��1���Һ� ��A_�@��+̍Z:�%у0���f����N����S�޻a
LLk��>��ą��ܵ�������F�xϡ��{���� (�>�k�����F6㭭3�Ɯ����|J~�%a�Q2��$H�E��w��-s��L
�X~8|
*0V.��d��:t�i���}F���S�6;?ygc��U�L�!���T�~��%�������!��M"�ݾz���P0r���U�؂�h�[Z�?e᰼4�Ʉ��J��,	h�4	T�򼀼��}P��5�A�jgl�K��VfmP��_Za�K�A��+95��t�=yA!��#�u(� G��I���^ν��wt�AD����ͅ�VK���?џ/�,r�D��t�=�L.�r7c@��Q���(Bv���g����v1�ڻ�)���?+��ϙ�?��Ң��
��uF��Kk�1����uĦ��+,da�d�J��t3�X_Z�w��W� �V1b>�A2k5�N���BFe��]�Z�/N��r.2�xr?1�F�+h��t�Uxך��ݽ����/�!i����ĢPL��0r!��.��+w�F�.��0�-�$PAg�ѧ�5Ś�^�`��4W�v|.l�l7�[�:�f�!SQ�����R�a� �@���)����j5��J�5B�'Ga�tJ�Qu2�YZsF�&5��dJ�q�N���w�#Y�]�d�<��������&�S��]�z�u�$x��@ú��TlqO���������4�<��l�����#*f��|�.Y�r�̪E��fI� W3�#	񇲆!׵	�ו���C��� �K��Q����7y���������y�E�z�7�kݠG,�V���C`Jf�|Y��~��2�-�ڨ���� ��\�_�fU���`P>�/)���E�e;�PJ3�[2�j}%:>�ఙ�Yo����*���-�2=�Z��k,2�A�t�'Ԙ,lap�{�C�1sG����ҼmA[}9p}�������M�=�My����[�D��Du��b��%��<�E� �[��I��t#^��U��0▇6�G��E=J]�5�V�a���7ς���\�-��W6�� 9���O@PT�ݳ��f�S�?+�,�}� J�fJ�0�`��i|O�y���(��u���sR�t�����a�kӪSԷt'�s!�$��6�t�w�ns�S����a4��m1k�m=������>��g����4���0�����*��>��O</�ֹ�z"z�&����Gc�j+��=��ߴ����A���Tr��0׿6��`S�%��0����K���4�g�����C�lvi�6��vI��>`�R7'��挊��.���������3s�".�3���Bς _����{f��缛�58��ЪB�6ܬs��mM!�ŀ��oR�3ɾzE�i'qM�m;���<W����r#"������tX,�?�2�[J%�3�/�Z	K��\���e)xx���Y�N������⋓��	�R�l�n���[`����P���nI��`trz�VsT
B��x��t��EO�'�9�6f��P̘^tD��%��z���"��V\2�-~|��rfe��i��H���l"�L��4�pR�^���������rV�kC�.m�@�3ĵ�� dF`ڗ��Ŷ2�my�e����+�N1�W�`q}�6vD�y#���֍gH% n���?�+����CI�+�g�F�26�e h�ׇ�"��� �_D6P�����c�Wid�Ǿ��N"�u�-~k%�}��w}ܳ V��Ϡ�mj�Tl��)�g�ӂ�	S���tC���x|I,���<���Rl�6�Km�ULZ7�� wǮzg�7��uT-��3���`��W�
��A��1/$�ƍ��σA����ڿ���Q�qU�J0+Jvl���x���z��Tm��.�-�:��20Jy?�5�)v5w6?�Z5Z��&�� �W��9��!�M��q�4���N�0h_��zl�`�Ǘ[0��\�OD��^��N(~��e�������T»Z� �xg�rB
��:rEU�/�x8'e����L�w��Z2��Wx���D�$y�z������޷��.x�s�w�:.���H���nׄ
�R���#�|.=�O?�,ɂ����t���.�����-
0�\�,���m^�VT�ȵ	d 8�>)�� &]�H7ä���~#�"K�H9?`���N_@�W�O�ǵ���%iP3�5}i�jy���|kb�� ����<���*&�"Nw�Ȃ~$�'xCE��߅�KO���?�Q^�=}}��it��l���@��^�E�фC���Zޅs�"�����W�����Pso���gj]�"�*���m�N�mec���xi��5�P�l$�&��ǡ�IC
(�w����'�_:�N��|�ADԋ�)+[̔���F�oD�
N%�֨A_����d�&6'���%Y$2�r�����*�$͎�S*��؇Z�@.�%�X�@�D||iX�-L��	�FIR~����9�p"<��erϼ���c���/ϓ ?��{,x����ܚX����y���I���E�l�P�ld�քXC9�� ��f{�]!�ss��ߋ݉�9��q&A�]�5$`�Ǐ!C6q))[����g�?�y��Q=Ag���� Ճ+vI�@Jq���3��<YhN-�lG�G�o��p����T�'��`o�\����!��p�:�6�!5�����8�Z;�'���VL��oFd� f<6���Շ�K��Rl��&*�K�f6B��o��8X��q���!
�тMA�+
��*�n���" �MpuJ_�h�����H��_ݵu�b������N�����݁�0�{t���A���.r`�pϵi��gRz墨��#R�����D՚I_�op�����	�U7��Mq,$�Е�1/9��-�� 7C�3G��HRCP`U@����7���hdi��<]�����.P�#��� ��$[��%����E�Y`|��\=2�᷽�G{��1�I�K�I�:����k#���p��V���w�!q��t��+8i5WD����	����Ů��IK>�)�X>8�nNH�7tb�C���[]�E����leX�S�k|E�dJ�(�Syn��rkn�ͩ��^�6��Yd���.��|����6Ӽ�<�=zw�g�7�?�@*�.����I��,����s�$QZ���N��m|�ڐY�`D* lmc��iǎ�0^�����zo���$��4��!>�:�ia���sה(T㠰�\|�������K}N�(��9ox����qJ�&��Ϻ5�.-��@�~�(���|��s�p����.�9���/�Y>$��b�w�ԉ�l�U~��%��G|����3?��7$��HO���e4���Fs &ݡ�f(W/{ X��^	�ޓ>t��g�2��(0kģ�t>�]U�t��!���rнBE�+_��C�Q��A��&@����刪�߽
�+�#K:L@{_JƵσVv��;�,�b�NQ�2�bz��#\��c�y�%�lq�+-��O�@iq4�֛�_(��lt!sS���G1A� A�C��&!�Ou���lJw�y��U��<�2�Y���Yϰ{�C��Mt�on��i��1�X��D�(l-S��M�c���N%�����"I�����ׅ5+����v�3-N�!(Ҳ��E��N�(o?P�
AQ�s�{��N�rm���?��<��Ṯ:�f�j)�z{<�����"&#��4����L�YS�6�U���=��|�/&�n���u{I8�.��_�T @B�i-�ˆH4��'�E�d�8�j��gW�^|W��,0�Մ��2S=�۵:�n���,.2��г{�����Rھ�H��CCJ�xǣ@@����j	qT�Ai�������b�3�&�e��oYMn�K��3M�_X!O<d�e��p�M��2�h�=t��v�k1a��}Z��B��ez;d�0re���{�7kU����u�
ݩ"�gxJ��7���'r�J�1�!]*ɘ��<T���1�Ũ���1�q��.�j��"���*���wmӃ�$�G8�z���s4�A��%�/� 1c2w�����K��%S�k�i�O�Y�	�
�!rV蒐_�i��HsJCJ�RNp�!��14�I�d��4�-u�[�X�e�"�	 ,U����1Y\}�P�l�����Z%�K�����j�1b �l�c8
��P N�A�х���U)�G��͕
�Z�$)�,}�_\p�Һ�;N�x:(�r9�o�����i4�\Ü�2�65n�C'0�Z-]̿�{n�(���\��MaX:�axM�c_rT��ĵ������� ��u��4�GE��'7���߶�FOt��s}Xx��ӓֵ��"���������|Ǧ#E��0�w��d�ө��
}��U\��MԱRd�cg��#c��R��y)��D=i�j����Ⱦ�cT���h�K���P(�%:zމ	�K�ǃt�L��g�^Ep�~���5%ׁ�H"������.��b%V�|(��+��nA�)1�k�5%��Sf$L�Kk�"�v�tw�m����+��I�`�f)��}K1+r[�M����c�6�Bc����H�����E��Z�]�L�CR����|(�pD�> ��[�!�ay�A��o�V}��T�"�0a���A���~����c�Jk���!P@X��qʭ�T�v�``WB���N�µ��B�kcZP��?��q1v5Db���O0Q��Bo]�����|q� ��?������Z�r*9�u�Hu��iR	&�;������ЪfpKO��s�ig�d�9xj���
�o4����b��hԛ_�h�}��2M�K�m�����5���ӯj��Zi��{©1��a���<�������רb�D�lk@W�[3�-�?2l�e�>�첦)��&us��:L��
���\:��gd,9�����}�]q	�Y;TY��bݜ&�� ����Cmm���ko�L�[BVnzã'?�6�L��ɏ�$)U�[�DIL��a\�o�2���9�3 ���ђ4�/��>����-m���~��V�m���S�_q9H+��'��ӷ��3��3L5�N1bc�}+�<p����g�A�JBG�m��,	����(a�0Z��֓�� �]1�EM�\p0%�|���N��A���w[�gU�al��?h��1��.�����Q^�@oޏη�l�6 �z�TK��x�d�3�')F�={
�y<��J>{X�ԏ���������*d�7�ڨF-�Рl0� )2҅���h'��J���ܔ@,k�}�(�ݾaܗ[�D�������q��L�.N����\��D��+:��~b����$��>"��%���+bD�5�ڗ,&�?d���c�$dD����
&8�\�޵<������
)1��Ѵ��l�nlR`���(����?f��&+<���+*�x�����r����*[��G
�s5N"�yAց�Z���
�8a��k���%V�LWӖ��?3 �����2t
�:����ƌ�H��TK?hhWY����ړXH���I�T�#Pwdco�IQ��I����K�KO����0c��`��q6�r��^`�����r��(�4%�������Ω��DՄ����+)�Xj����]B7 Qy[�	 6�5�;KI�s1?���Gy�!�{��J��^rbxJ�ql)�W- �>��vu�y݉):*�y	"�R��,	�U �s��鶗֎u���U�Y��S/rxrѷ��9�*�/}]����R�k9����f]D�\�T>��50�!E�/��+���w�rM5�2\B?�D��yd�Z
��rm��m��l����,|���W�E�:w���n�Z���C��ق�J��,��$#[=����3����tu�2;tX-����x�R	�V�̬<�����p>��,®�9�)��2�P��`&U	��Qv�iϘ]2$����>*����|x��"���'�B�M��2�&���!�B �r*aMB��l�{��x�L��B5��+6�m¦M�4=]�+�Ub��K1��I��ؼK��5͒jί\��0�����r�,T�GCUbX�<5��b�84$ӆ�Z*��'�*z���EU���8��<HP��ȋL�F��®�h\T�R��WB����'�m���m�A��r� �H1�����^au/��ڷ.>���-Jn�H�
�С�ٴ.����y��HD=V2�H����b��f�<��R�G{I������k =x�-�d����j��(�C&�h�c�S��&e6B!��IPV��B�ÿgw��T`р��uv��2͙���ѿN��J����� D=x�ߙ����{����KJg�y%
�ա����c�wW��tI �h���"��	��������*���t'��^ k���ί\G=-� ����?�N��	�Py����� ��4���t=����u�k��sϘa���މubm1(�ŘL��؂�>H�&������*D���T��AZ�cmM�N��*����������>Y%��2���Ɨ�kHs��u+9�,�d��'�%��f���u��H=�\�ޭ�����A&��@hd���Oi�)�x�斵����Nǹ|�Q�l�������������-��~w��u-������~*�������,ɹ�>*�O��/���EA�h�.��4���&[�	�YBSK ���3Ц�z������z5��k@o��9#�������E��G	H�\(�/��ص��%��ڣ�I��gU�p���G�΃�^�e2�����������x�d1�jW/\���	������93�nQ�,��}�u�ً�W���8��fdʨ�&��'�tJ����L�6��F��]�>ؐ�u!k5""���s�s������8 �7��1�*{����ͻ�7]_�5�;\��D̂,�'|>T�z���?���sƔ��ǅ> ����i�:�����̈B��wG�a��sg��m��PR�����G�?�^�a-|���T�v<g��Q����F�dfZ�7C����SO��;�1��8@n����Ư:��J>U�V7�㘓�q��	,�����`0�]"2���Fm�+�� �+����L@�}шU��;#;f��Cx�Ξ�D��p7�=�'1a[H"\���:�]�샶JIQ��w}���s����>����W�=x���GQ���k�8{Z�[���^�%����W?Y��~l	h��b₰��H{�v>]�u�̵���?�r�wh�R�9:
-���,�.7��Au����n����o������wYA�}�¥@S��C2���wV���֔��gNB����7��QN���"�?�b��k�w*����	2�<	sz�!1�]�~��I2�w!8��͇���7�s��s�{�����l���kGڍf��!���	\�e����+�9Թ����C�XL=�4��=����|�&s}���.�)�$��6 GV^�뫰��m�w\�@�:���N�^CY����aLsB�fWyⱝ��1ej������U�
-����&��*�9�����|%��������-��"���6b慤oÚ�ݰ>�p�f�٥��Ǧ�B�Q�pZ�>��K��sН��s��̯�����
 t|��ߎ�)"�~�-��u9����k5vL�'�:b���c���(�e�_��8���^�b���������Q���U�  ���P�O�7�C8W��Z�st��~;$�3.ѝ/���:��<���4����!yD�V��©�����W��o��ш���x�L�L��f�ʈ��+�|B<�Du ���&�ƚ&.d���� �2JE���^E��ѻ�=�f_]O�X��f��D� ��j�)H)�������S����'�����)��"�mB�il ���uNsի������d=�����̡���^�K�
LL��NE�Z_!����g�����i��gUu�HR	�D+i���Ƭo���U!~/n�4Ͷa
G�2N/���}�H�2z/�p�F{2+\]�X��F�f�I�E�-���(B�������l�YW�䌎�P#�9�C��! �4�qј���K��:�g�Sf��d�͛�Q���zf7Ȩ�J���2v)�"P����L@�5j��eE�v����V z4�YdJ�21Г�%�ٰg�j�+*&�O�(0Ü��-a/�Gu3��m�sȌ��2̃�4q_��/~�֚6���@���pQ2�{�/|\��-�o�K�D䵃��{6/Ϭ�������4�Qu����y�yc�I�����`<��{��f/���j f�s���t���FN���R�|l1�A��2\j~�.^F��/k�x��a�����6�(�Qx~��Q��ky�p�,�3<F�o#�Nl�aո�������̼�%|��<E�¾>�R��A��	���U"��4���$]�{��o?�{J#��'+�U�Z�^EG����Q���E���ٺq���d�_��v~�}����C���9�����۷�u1��H�������D	a�`�R�̹��U�,yzJ���q�r��,	�=�B�b)t��:��]�FS�I]T�ʠ��:�UN�ס�ʌ5�V`�P�s�k�0os�{��m�9u�ϯ�S?W�$M8��X�O��;K���|�o]���1r�K�F��NZ�'�-X�E��`���˦o �?�q��i}8�ؽe���]>^��㸭�a~��GN;i@BY3ݧ�
�׀j����w�˜~�W��?nz[T_�%�X���&i�:��DZ��2�|k�E�{Ơ�c2�[�(�4:���4`Y��,��ƞ�X+T(*n����Q������}��tE§���P(K�Chz�O��o��k���8~�'��7���x ˦uP����"�����gV�|���v�rEG���C���*��i��dc��-B,�9�k�T/T��O�A��~	���8Ў1�,"�8g��f8�%Kx�k���Ne=>�fT=��!�"�c����i� BVLa)�I�?<=El�=;��5���b]|s�ߒ�A����b�*]�ټ����qS~�D�9��٢=��q�I���7�_O�B�W{����}��@�њ��F*���_ڧ��?M����X�GD׺w�@fq�^3E�����qX>���bV�-��H�NCx`l�|��8�p2='�7�/�=��� $�[�T��.$�����(�UbU^��{;�j���l�S��:oX���W�-u0�Ɏ(�L��u�X�*Y���M���oT���E�R��hK� ��P�Xc�Ǧ󨌊�z�T�6���Tl�����;�m�K{`���$��${�[J+�2ܔ!��Q`����������"���c/�����6W&b!�tw��}`9/x��B�=�s���ߏ����=I�+!��F?��	���ʘ����3E/�S��`IĠ����n�p�H��q��ڃ��Er>��wO?��������)�j%)�Y7@�[�G��������E�^�S�O-N(����f����nW:1�Rb�Z��Ƥ4������w�����z��ud��8e_�C�)��"Fy��E?9��BQW�x�#k6s�<�I����x������T4�6E&O\6��0.�'G�������g�\�����M�;��1��n��V��g�î�K��Q@j�A<�Bds\�P�	x�2�%\��>�������Y�rJ��9�vJ���LX�YǷ�p��8�T�Hץ�b�a����p��ш�=Dgb��	�Q�o��`}l��[�A��]Z
���.���ЎK�奺}���T����9M<n��Z�azI��lv45Kp�7V�����<���D��}�v��*�Q)�hG��뿯���+`sK�rA���/��.#:�S!1> $�m�PU�>O���S,n1�m&뺄}�o=E]d_8{4ѭ�Va1�B~�x���.����5��pE�JL�lF�H�w��1b��N��j�pU5e�0��a�`L�t�N]�s�/I,��M�4j�7���������g��f�/��Z:���h�b�t� �9����jC��H�:�3��x-z-�E{� VY}�c�Ɂ:�GƎ�^��Q�6��q�^��]H�{#��7o���Q6_?9I�5�!��O����h���nu���y�e9&(�s��2��e
�?��C���wЮ�{Ԑ�4�aq�'��M2�N��g������l�Z]�#QXV�\��|r&?��lm#��UƉ�S�m1Dᗸ����C �}2t��0"C��\�a�y�aQs��O"h)U�,�nP�Fr��n�
=�:n?��9��8-�tQ=n�9���^ٵ��zEF��+^�E�'$�06���:�~���b+7Y@.�3G��	�V? �}+G7�M�%I,\��4*W�Ά2�'��
t6��uê��c�E�n��W�f���(�!�j��dJ�rc�����'lV$��YZ�=\7�E�dɲ�)'�$��Ȁ�ˌ���ϟ&Ӹ*�ːR�B_]"/�0�������6�>��9��o �l �9 �J�
Gl�|�>9s
����wK�Ob�q}>�N)�q�/7SGi|�	�=��L�|�������L\��8�9ӄ����eG���KWmg������5܄��c����%��q{�kO_P1=�Sdؖ�/\��2P�Һ:.�b��W'�ݖ�/I>��:*���zE�u����'W�|�����Y�b_RO�C�ܮv����Wo���$re��/Ԉ|\14�]����jm�4һ���1(�g�@j���/a����J��G�����8&� WlSB���k|$ c�CO�LlfO[��Q-��b��}�^27�L��r)�xr��rY��?�\y2�0�[�3S�����S!��_*�V�ok�7G�B��N�\�һ3��Z�)6!����(�-�H�L��O�(F�+NR�1	y#Xf�ր[؍iyT<;q�G���ЀҴ��q��S9z�!�D���D�di��d��y�fi��T�2��2�)u$�l���)!��r�os���^ T����zN����g�u},�t���7�l�y���#SID�p��e[+aj�a�Ut�(�Y~��~���~d��Y����N�`�u�'�"q��t�1����Á;���.��`������/�!u�*D�*��`�0.%9�J\�>�lkq���b�j^Kґ�W�aLr�p���W�/�p�te�V�X�,�2�柇D���?$��nwO��-��mз��h%�B>�Ȳ>��(3���;2�f�W�����w ��	(ࠇ'��]�����v��j�m�:,b�f&�V'�xHu����M2y���\��f��	"~�@��W�-���y�ԧ� ��Ui}xE/f�l��>JT�F�@��qT��l-�:����W�g(q6�*���񌊀ry�|�*Q}�A���~��̠#���Sk������f�
=�R�ֵ��9�� �9��n�X��?��?P2�ד�gr~Z��)M<H�X��!o���pΛ� �W��������Z@�m�ب�������f��I�ƃґ䤞FӧW���e[1v�����(��R������޷DW�������91�I?�H$ �?�L��ڣL�K j'�5�O�F�����[��CXH�� �.��J�Ź�l�|���ӜϢrrFB�S�M������Ք;���O��
����'Ą �N5�]��h/J����X��������/Z����ĵ�6hK��vQeж���k�y،�Xo���K�����*)dF�Z���T��o�,S$�GK�*�l�%>>�_��^9!l��}6��qM~��=�cg|���p$n�Z4X���l���k�qIK�C�]9�<����Y�;]��̀��=������Q�ӕ����:'��X���B�5��C,;��@*�6+̰7�3�u�����@������'�D�:=�(��E��sب��Y�ƿ̋���S�7��J��b3��1,��=�<�X��v�%y*�h�`������ȕZ.�!���EDEj�[ܘ�q����٘��|K2�w%�Z��Z��4\�)�A��}/FZK�=B�
b��@�A��OI<mP��53 ���[~�9=T,x[)bL`}�
���9Ҿ+!�
j$s�z����ch<�:���)��$�� MeK8��Fa Nދ���)�sP,X#"9l`8��-}F�0��n�pu�\ci�i���b�?(ר�~��H�����J̗U$�a����m5(������T���O�yc��Eds�h�͵n©���|7�s�V�BXF����$x���h��JZ�#�{0Z�?�8��@���6/���]�*�\M�'�:�"k<Q�/����� 
��V�i`�M8"U�K��%kz�bn~�Æ�;��+Z�Y�ˑ!�v��y��I[���5O35"�����;�m괱��	V�2�nރDU���q��}����[P8r�v�fV���w��]�:R�N�d�q�!�4�y5M1�D��̑B<~�pmu���~�=&&���`b�'�.��"���I~��5P�C��[���w+��j4߽g����Zj���#vԤ�~��;Jez�o���Ah��5��@��ϩ�q@�0:OSKLƍ����ǫ�H������O*�[ě��V[P�Ս����@�/W�3��C38�Ԧ�J�,���p���p�]P�
�9�$M��\�[��K���L�;8�2���_�5ai0�/%s>Q�`y5�(���\��M�Z�W@v^+�u^=��>'�O��ϣ��l��q���hd�mQ��d�H��Û�F�67���mԂe���/�N��ʸ�E���}��\������dU�)�����-�����d�^�hċ=�`.Q�H8& ;�6�o���%�R��)�x	U�G$#���-"���Sr��o����ϱJkBS[�n�����;�{F�`�{��Z)� ��M��lGg��X�h@�S���&�T ~�� ��	(߮�q�񀬋�\�����̺���
<����[�!r	�t(��T��l����u�pF���y^IO�Fx�{P����0r���H�Lk;�PY���S?�p�JG��hPP���L|�=�4��'��w� 4�6��[�T�^D.�k�������P�ta���7>�9ct:ΜK��g"[�Uo�$pSkSuF��$����`�z�I�A4�$}+S�?R��9� ` c�����!J�B���tՌ*@��Y�2�����=���b�s�^ex�r�2j��=�\@��#�D��@]��w�%��(,��82����N²�*J�qƸ�/
hM�RVZN�F5aY_l�W�?�#��?�+�G������M�%���~+��%��@)y�������J�{��0Η�P"��J���\�����>�?=K�G�bp,�Wa�̭4L����Y�e����m0�L��j�l)餼�I,��*H�?��tC��ra�m#Ƒqb���!�6;���w�������G7b}�1��~����\4�Pc[�	��|a:�J�����dB���}<+F���؞g ���(d}����[�����)z��9k��w*�6�2�[e�<�ꀡX���{��[!ly�/����U�'�K�]d� 2��)J��V�b����$o;�?k��]�ɠB�!at՘ Cs|���P�<ޯ\ͤ.ܲE�&�&�]]3b!���ۼm���CI�^z!]�&4��/�9���fy�ίh3�ݚ�x�ͽ���8�t�bʊz2���}%&���E�A������4NH�3�.��0ɳ�[kc�>�F�u��d�詏�.p���	N�����6tT�V�)q�#�|����&��R��S���-޴Խ~�\
�e��Fo�(e�W�ꊚ4T���F�2x;4���pjk5��a� ?UR��!M5�L����jy�y�F�(������4����=X��\��h��(:�`;$&"<5'��ga������H��U��l3�e�ThI�ES,- ��1��ќ�|�k��F��7iC;���$���)��Dl+�62j��M>�-�JmƱ��i|G�y��`3��eŬmk>����˪��г�B�(��d*Z"��T���Jg<�NiL���K�K�6T>"���=#g�������,�X�M>���-_�x;��X��6�vx��b3�jc�-��<_�?wՐ!F.Ϯq�s��<aL��kZ�'����n���y=;��tj*�C���>�R�j�D�:W���Q̸h�N8�_)?z1�>Wbz�OSv�ZK�Ik۴�% ,"�����Q��k�|�d�tНf�������~�L[b�g��b�F���Zm������ۆ/�O/j�MZ�F��	_��M��or=-���uR}3���L�0�EI�FLJ`2����OJL����o
ł4�~�5i����i<'�}�~{z���`ZOSy1�B<cc-�l�`����&N�-���q�R�f�gq��3��2`Y#d�ík���������1�Xzk���G6�d��$���\^

��y1�|"mR�I*�V7^�<�Λ��#%I&�Zfz4ʲߌ�)ee��o��x��'0N���K��mI'ĳ ���,���L׈Yj!�����`�r;����h�3dRI�g[�ߴTb�iL�A��2F�v�_[�QH7PS��I�TT��Ȳ_v)��z�ܠ�Z-7�����:%��콸G���$�j9 Mlv���b�e�f)�xh�k ��'~�\�AC��z�Ǐ>���GT���3���x����l'��7_A�zj�$�n�SN�(�ZP3E�Y: ���S�[R��ڈU�ye�Z�i"-�<"	��ϒpA"?;)�~�qi�9��o�Q�Ǖ�R����Pk�uw�8��%t���iڏ~�2�����ڥK����WZl]p�}_���K�mm�d��)>&��N[�&�1\s��;ʉ��_�x���9�K@���#�7�L�b4��$�=�d���S��Q�Ο%�S8pS�4����tםX�3d�&Z��������>�|��>���C�4���I�񷞑P���y�c˛��$�Ɍ�����Aq��J]&�%�}Q1Y\�T9�d������G��i%�jd��G3�GKM��̣V;��4'UM�x_����@f�w#����Gޗe��G�Rj���Ū+�^}�ļ�64Ln�����5u��� �n܏!԰�a-4�>͖l �{����-�T�W�CMʫe
wr'K.>jdwK[���w6���rbIȪ�tț�;\n�J ��ċ(J�(M�C��Z�)ϺVz�Qey���A���o�9<�m��q�E�G�k��7J��0��Y�F���rؔi\�Ho)�Il�kd�Kñ�P�Dy0���)DW�~�����sXжH�>Q�s�S�{'�3��h0��r*u�j&��l����/;�8ZEe�+��2?�94c���C�^ף��}T3�Cyi���O���a��᷊�����< ��"���;|ݼ�_���\_݈���)��롘��y���66��L�኱{�N`��G`��d�.��btZ"��3�u.�|�R�еCe1N�&��9�P�=,��=�.��n(owط�H�wx��ؤ��x�G}��]�*'G�BC��
����tD}Ԉ0��1pW�
/��Y���*�߅��^�Qܚ�Y�L-%d�R
�k�k��l����Wz(���܉M�{�z���]���i�"���Qc�:5ɭ��7e/p��� � E�[�nt1!�F�;��ȧ���D�ߊx̜����Tl�v�$�^8t�����p�sh��r_��R��	A{���ZV��MC��E�]�FЧ���+(���t}	2F��rr��������s87������3����SUf�fl������kfߠ|���u��#��!t�oG�~����"���!���v���_#�w�����&yHȋ��'�	��R�Gi�wbs���K�F��. i���Z&�����1�����K}wb����f'����?F�A*��X�����U�Q�����%�J�LQj�4�`��̌IC�4��b��2'��g�:y�K#7�s��%��#�#���)��͆_�t{N� �u��p�N������<�m���߳5Ifo ƌ=m-�3�V8�����#��e5���������
q��-�JNb!�m�z�"�+��T,�d���au�������ã���ip�cf���=ŏg�=��z�$��$=��DNd*���@�Ȳ�21��?̀Z���	ʴ\��\�<c'�A�\�
p�7�ўR,��ӿ �<���-�;��X���Ѱ��m��\G�~]h�ã$!&_V�����$(<�W�N�{U؟5�z=3*vv<���NQ��L�[ft�7�6�����OI�(���,O��w{�K���պ*�O��B����G���2]�|l�[]�$X�?�RbW{���igkS���:1������oI|]9�"줂fE2�LSK����&� �t�CTt'�Q� �cD���	~�����Gˁ &5��=�{@�QHB�W�V��iW���F�D=y�7%
���Ģ�d �{1!�E�r��Q�	b�5���լ���O���MQŰ%j�3	��_��4n��5����1Ng]/K���r�=��
<&s��"}�a�\��L^|�α�ͬu�&anRwjҺ�g�@cP
�Z�r��p�W�˷h�a�0�/?�����i��/)�� ����a��n3�S4N����n���J���]�?t�}����� t��1�a-���pE�����H���I�S���ُ��wW��v�p�Q��X�(Z��.]g���>d���fr�d�7�;�Y߮k{�,o�?�r�Zs���-��P����ocDQ� �4`�HQ����	�C�`T�Ƞ>�*�nN��}!��'�t`���:�6�,�<w���{����X��Z��ԜbT!8Z�OYݙ���?����&��A�q�g�#ȴ'�S��d7,34}߭�X�ҭN�����A5��ƕ�?�&9�:�͏�b�R���?+$6�� 7I**F+)�)	d��̘2Jă,w�Q��5L�k$�Ys�/�v�"7pQK���B�'dݔ���Q$P��G �I��Ҵ�3Je�Gbn��?�r��f|T�t���;/X����M�>�E�+c����e��N�Ӿ�vpqƵ�Vu�f>N��lR���v�gD$zv��&n��x�1V��i�;@�.*:�I��l�Y3�j��[���C$ ��Y&.�;d��+rܗG&�O5y�=��B�Y����
s�42x��ϰ#q�!��%���1�D��4"�:\�.<)�4�;k_Ho`}ȥN�l�[ɮ>�XW�,��v	ZSB�Ĝ�� =����3��,�ը(��a*�O9��Y����٨*(G����U{��W�(�~|O�>�tK*����ekw���Ƈ��
��\(ڪa0;5L�e �˽����������/�����ȸ*8�ݠ�հ��9��Tr�˔I���E����)/ ؋��w�,&ɤ@蟁�qŅܪX��M�����NMmG���xHW&��B���|q.C��aHt����ձ��s��`����$^�#'QF;t`��܄�+#Fטz�{b��t0Vx�M��n� e8��8�M]�)�|C	A4��xGqʆm�ԚJO��,�0<Mu��&<� 효*��R�i���&�3����������4v�w@�(�"�(A|�Zx��k�m��|�r��N�;��"�t��x����(�S���r6$�o	f����E��ҳ�;ړ8y�?�7`�.:�i����H�=G|�����Jv��3�ڬ����^X����y�}�A��Y)�.'&͉k��*��zZǸ��袃=G�@d�!� �7�-�ܻY���|Tʲ-/͙����D�{�{��DȮ��Qs�Q�6�� f��:��T;���Z����$�v��@}�f�'����'�oo�R�p�%�ч���5�+�>�l�)_7k�C���>�(��'O	.��$�l���M�ռ�e":KU����&J��dNg���nIXI�8�>��4)�)�p���ՓiLY��y��Q��=��'�~������p_�j���\˕a��a�]ٚ�{��Z��Fx�m'�BI���풢����Y0�mӊ?�34��M�Y�9�g��9 O�v��Ƹ[� ���r,:�m��qt��c\}�B��uE���W7�f�㫯@�0���l��f5��>��/����E�����g�7?�`�L�F��5��#�ͨ=�=l	��B	 U^���f	V��i{c'dR��Z�3t�� M(�75�	�zw����Vjmq_.H5��9�5�B���͒G4o�ʃ��,��(�>!W�g-�y�h��r���V���gá�|0���z�'�d���g���zt��P�74`+f���C���fE�p�A��Ë�e8:u�Fm�]ڊ�Vi��n�&G�fH�E�;�˭V2�+�>}�P�p$��񺻖�*MlL0�I��Vvn��2_oTY8b]��x��o\[���߁�}M�FrB�١��~R���<3��r�j���p&_)�g����hi�0�P�ii2�u���̱��[aX��=խf�;&�.볭��i	|0�}��ۈHbW%���!R?�:��u_o1e@�h �L6�X�8���cs���0���A\�0���������abqO0��|��d�0��%c�p���LA�x�ʭ�����5�}���y��m�}�?�7�$�V���T;��!��R!�9�o 3�K;�'�$Ұ�K������h��`m��&+��w���QF�o�"p�ړ�.��a �n���j�:�#�9iڱ ��"\E=��_���7�����E^X�V�K X⿀Քa��a�T��V�Y5��bV���ȸ���.����Ft��������Z��[i�B�,Rro������9@�՝���?���=�m�s�J��&����!>X���4Oi�~d]�qH:���8��Jd� �$�� ��SVaj}��F?�[��+�~�&�=F�/^¹��0$u��6�;xKj&Q~��7��?��
t��� J�d7d�a����=ͺ12���tp<\m���\Ǣ��e��B���Us�����ݟw��j һ��ya���j���g*�D��x��.��;��mN�����G �؁ �!E6��nr�g�Ԭ�4�!��Y��I�r�u�w4m)�2�>(�6v��?�&����:���BJ���5y�J�|�N�K�S�a�'P�r�#e�GMݑ����La�`�,y�/|��9�͢S=:�c:��j�|B�Ď��-���+E:c{}`�<¢���6B�Q]*��q�Xz�;<���aku���8�E��0"Q>�Dn��Vyk�m��j�"g �	�@���B�=��F^X�[۰u��
$�+�֦c)�q�s��CK�k�og�G�Iε�J���2іO@捦���\kIh�FI��e����,?���#/a�I6zI�h�^V�O�O�E��JY��>v��:��O�zR�M*ߊ3���Y����BQp��ʈЍ��iK�;' ����k��V'A�~뇢�ۓf�3�V���S���e6��,w��cq��⹛d�m�����)_t���k�B�G��,��:ɮ�z����s�%޵�I��K;<k����2�f��xI��2�A�b(+y�G��V�G"pGLgݿY3�����:N,����,S0�Gi#^@x:�{JY%�xb�	�����x����3BT�yT��Bd����ƃ��S�G�n�;c��q�t��!1��E#ɸ)bW�7�"���1��J��l	��8���tHR�<�N�H��Zpa�D��d@�v����m�j��JΘ���Ү:l!�=��/
�bB��lz���xdC�y6�'̀�P�0mQ0�-�����7��7����V��2�R1K@_�LA�D�k�^!6sIQ�A��"I%�엟^c�Rؤ����� o�]�ާ�h鞍B�*�4~W�����r�&���ʊ��K��=��u�--��y�@��+~_��>��=r�@Mo!M��3((/'M`��C5�%YI<�yq�7[h�17X��� ��8li��P��f8A���	��;+���J�xԷ�Ӱ�x���������}p(�Qo�7Cv�S]c^:���`.��3	_��ЁZ����Pu�r�� 7s����$�\b�\.��=�x�ʖ��#g!��c�ug�8�(�`��*��,�7�L�+�!�i�����6�&'�Ex+kLt�E���Y�������f5�`_�:Y�E�I^`��p�C|w�$�q�v���De��-aO{���kȫ�o��銝��w40���!G��h8�R<Q�9��~�^R�H����(�=���\| XW?�v�`����u�d#�0bA0����Z�<���!Y�+%.#ŧ�<cUh��}���mgP2q.�^I�F�M��ȕ� ��}�Yn�=�t��k���K��f�K��~:�ߞ��jPV�
���Xn�/�?���I�b����BR�=EGf��Rd��	�� �E%�N�]��pE7ho��9+q��~�ܪJ�/��
���Tg� Mu�}�~�b���x�
�g�>��)�+�1 8��� 5b���j���l�9+<�`�N�8�(��D�i��m^�b��"*���RՏ�ĉ��B��E_��=P�P	����I�Zmۆ���t��i��_�� a%O`H�L�__\ca\����L�q��BRUq��j���_N:�hb�2�&��D��# ��V�>W���P��~��=�e���ZT(jZ-�~�艊�y��&��ݎB4���N�`غ���X��Z�>3 mSվV�q@#_�B$�;�^dZC=�c0��$�ʂ�sh`#;�2C2�ѵ������01�����rk��}��X9�����_�^�){��}���93��F�!gO~
]���!Yw��C��&��}��;�20�p@�h-��K+V%LE���N�T|�Ω�1	�]^��;�g����F0�A�2C�z��vp����#H�8�-GZ�Q:�%Ȓx)[�e�=��:�A�G����&���ʒ�(g���%�SpG<�׊s�/t��xpb�"|�$8����"���i�9X	&+��nkz$Z؍��d�W����e�F5�?hU"Z�5�DI��YD{E9���=�{��q�nV%�O5��p��-JK\�dfy���!�x�D�CZ���<ay�Z}��BT�7-�Y=Xc�>*�����w�燎�΢�o��>ş��Q!;�V9%��ڎ�ɖ�ס�z��E#j[C�O�e<h��5MTyN�u?l�՛X3�ّ�����+���AS�v���J�����2���K��Ɇ��|�;�ƿ 0~nb-d���K����L�v��d����`Q�c �U+���.�q�f%��K�B�C��Ʀ`���p��%JY�1��#�"�K��9�顤�&�s��J��uR���#����WW2�oh�DLH7ѽ�����Z����r��Rti&��U�G�c��ަ�䮨���8Z��=&�$�wN��V�v�Bǡ�|�Vv��<���y�	�D<�pԭ�_9 ��4�Ex�e_�^Ƞ� x�!Ue�n�*�)6u*X0�XN2z��g7��`�6elk�;�]tB��mw�Q0�g@��} ���~�('u�,�-k��h��l�t\��i��U�������H��},��ʋ��F��ԙ����C��#v6ٔT!�d���K��E}S���=��@�=Xܠ}�i	�!cc��\�A���x6׎�Ͽ�SFSo�`�
�.��3��iֲ���H�>V���}Z黳M[dܛPoc�P��o��2���fB='��o�S�\��N��c�CX.�W���:��b?+��ؿV���2a��k�r4H�:������M����P ̅���s.��U�#�:�{��Ԝ���F�y%?��~�-АT�&��<���j��"#l~��������9��Z@�s��R#y�F���\Ԩ�U7����Å���G�����m7:Y�U�)���_$�8(w�N�[]�����ѓ�Z+Sۄ�3:�{�<�k�����gp)�� �B��X7�k�¯7	��%�Q�K�K����zN=]�>�}E�oHt���Q��Z�16`~���u�9Ă����צ�?�`G�
�4�h&��78�8A<^�e����!�"�}�d[�R�ͅ4��C�C����\��yzN� �2����LDD��/�޶��a���������Rj�����I�o�k_�����pƭ��
���<��aA�G�q	�% �t�����;�@^�`\QM
�7Dp���+��5�7t4�tP��\�\{�'S����w���t2ۯ����8���oٝ�t������no�[��'	w��AS���vt�Wlnu;5�X�U󉅸�@������ꔑ�FӔZ��9'�bV�l�'�6Q���8#�s��QE�3�����M��9;u�l�E��fsoD�m��|����ZV����.E�g*X
.�.̟ lW��5Wk콂�s���E{���X�.�m@Wk�L�AH���0�C0�,�6�{}b�x����Z��d�ɣS(�0�~-���T��'�v�H4O���8�<^1�(�@�'���	��%)V>�Ʒ�� o���V{�Q��A5���1��!�6���u2�Yx~�{L��@����s�VR:�)�"]�mP�G��"���zr���\�M�2�4�a�&��42YZf����i�)��ݬ�-��[�Ρ�I���BUHDG�����o��g�%y��I]�b�������2��jg����[`����/�/j��<ݐ<;����
�)���A^1�E�l���LD��k��+��ۺ���O�R�(
�N���{�I��`h2�J�]Q(CS�]�g~e��<�4ZTPs��⾊B�\�Z���k��1�Cz6��,����5�kU�"<���o���s�fq�Z5��C!g�	��O<�o�טK35궱��dGUZu�����n�%�
��:	�»v�=Iָ_�"㞉�����!/?@��AD&�.���o��U��F�E�B�vWo|#kz	��e���V�!$G�թ#٦3���}��J'�S;��7��?G�j��_�n׃�69���C����Z�X��E�z(7XQ��-he��#t"�4U,x���Z6��Q��J\Z�W��ܞ���)�IR�DM���IQ�<ѿ9"���c������o5S���e��J�ce�Ϫ��ˍT�$�/{�g��x#rX��c��{|���m�M�xO��Η�R<�4���ً[�| �6'�����
����
��]��	�L/�T���>�:��zb���Mz8��H���}滁��)A�C�n3.�'����*R��737��~��ĕ&gہ�D�]�Q	�GX���(_ν?��9���01�����Xab-���4-��& ��;�
�f
��R�Q�)�*�K�(�WO@��?|�$�_F|�n5�7O
�/�o�%4�R��G�(e�������j�Y�gUEUwa�KŦ[�����3�w=S�Պ��h�D8w�Q{�)H��:Z�Z����)���o�Ÿ� �-j���L�V�tĦ
ܾ4j:|�v��((��{���t���{j�:8�s�1���x��+���yA���(��r����-U�Y� �d�;��� �g�C��ƣ�g�h�<��Z�M�q-��_o�����Vg��Sijg����6?h��U�6/�6��~m��}R���Y/퇯�}&�g#,+���m�̃`����:� �b՘ � '�U6]3QO�V*��˾�!���M�#�*��3��1%p\洑��Qq��:�Hb=;f���J�=w�u�u��xq���,��?D�k?�`�q�m�(��f����C��چ[�c*7z	�Y�F4Q��|v�Y)e/2� RlзY"��e3��t@�l>��
w�<@8O�{cEPĎ���KK?���;�E��=���0��� g!c�G�}$�[�]8"�ݍt�5�r2�`�ొ�����9����X�ec������p��=�ty I�h.F��q2��\P�H7���d��8`}���G�v�O�2Շ��"bթ�7��j�1�әm�)��R�O�L�G���^����	��'�D��}�Eῐ�ʿ����"bŷ�Q���`o�_ѫ0�¥c����bZs�l�S�+ە�s�i׋�@bοg���Ř��YV�c�Q��U�����o����"��(�������&I�t[>[�Й���Y[Nb|�Mˮ�lT�D�����V��q��	K�]�l�h�1x�$�d�'�~ۥ�����y�d�~J�ҧ㶤�n6F��3=�����z�v)Oe�JD�H�'9 �P��P����*[7/�������Glz��,y��YwA��0��|I��f���@�b�2��b���_W-x��^�K�+ɸn�T��?�^�Q��.Aa��fκ��}<?�Y���>E��t��� x�e�(��CP`���tq���#��,��	a��ezRܙ�� u~�c�[�Y�w���U��$_����̞�Γ򹖞EW�~��m2�s:���)���p���.�r��aH������`���eӱ��3�>��fC=���@��G͑Vݞ��9.�70bVK>�#����z�n���UOE��1�Έ(��̟���v&�I�ǐf��1:��V��J"Ll�M�|P�[W8t4�Sܝ�{�
�{话�U��T�<�|1';(�@xI����L�j��d��D�|~�'"L����S��l���d7���,�u���ڂ�%z��Qޝ+s!1��,JT�#�_Q��v?i�[`#�OK��T�/�=��)�V	O�z���S#UG+�}�&�P/��'c�s�N#��H^
����0G�Qf{(N/�E�{ZJ���'�+��8��zx��e%r,�esN�0{���@��x�����)Nf�䏃q���5��P��
��R���s� �/��2ɄExKB��}��9Y�*h3�vY��8��A���]抡�)��n�4��e0��c5/>W�Y��g��*6�2tЦ���y��#vv_(��E9l�:��6P�	X���f��|�H��i��עɲ�"��eri����c�,���)H\�Be��0r���1��~�e��Mc�Z�{�Nh�z�W �q���ɶɐuUb��#��p!e��>�{�~�d�)Z�����2�L�U&��ak�@��z d�֊
|�L�r}���䥉�E��dQ����e]�X���k�=�u���j:�yo�����ҨZ/��K1�-S�" �C��m��O*�'�"Y�b^;�m�C���SezP*\.|�]k&����['�JT�Af�۬�1�B���I�ƻ�ђs{ES�ֹ�^"���
��W*��vha�1;ƗL^��Z��0Sд1ba����{"<��B�]�/�y�K�l�PLeJ��/��"�\�B�p��Ҝ�C����K�EH�@ؖ�-x��6&��Z�ܬY�jd#h��Vƾpvy���/o{R!^�PL"���d����mN�v�/<�\Ae�b�)��w�f㷅�ZDv`�(l��e�"���p�W�N��f��-�TG��0S/�	��ʌ�m��+2}���Ӡ��$�u��x�!yu��B�J(s��L+]S!	���#���6���U��_��	�@+�衍fK�'��̝k���j��HJTdh�F�M��G]��n�:�o��/,�C!�A�N��[Ogc	2p���]��z�Tb}ܜ�&U���ž��_g4���<lM��]=A.���!X%��jҘ_��(f���P'�J�����N[{4��c*ӝh
�k�:i�k��5}�܇��nƼ�p\²6 4X_aC�[z���̣������M����2��Yy͘������۶��A�FEWM0�/��ŕ���b��Y.�x����12�IZ�����l�;�].d��Z��ǦmA�ުI���s�uo��2}��m�9Ϝ��/��Ŵ��Z���{�#��K��wH�r9�$�@���_�4Ƚ� 8�[)6����[{�)=U����_�O���7�����,/�b}��b��|$��Iug��.y8�w{��Rz#��d���:�>��܉�8sB
ڈ����TG��A��c��t����H%J�i2{�c�f�"�Ц�[s�����Q��[�0��r2ǻ�+֠Hk�����]6���Aaɘ�H�=��}���(���CCⅶl��ez�0e��v���.��7I���@��ס�]	�s!|n�xo�H��}Ȍ�]WV�{'����ˁ�i�K������F`��-h�]��ֱm��-��@K �� ���5�&xTSM����ܮ[~�sQ�6��|m��3�6s{�ޑ�����ՙ����Kfy�mI#i���WxI��U��8JP��O�H"�B�w��,3�G����`�P��bO|Fm��e&n�r�' |��E{�<��o����EΜ�+��;�@�H	�Q��+%�>
f]/�l蛘�f!�޺�L�����B�*�H�ܣ�䫢^�)��g�`�$�;�sN��ܱ#��jh�C
?�x�<,�\ξ����B�P/2T���[[t}�M���K�U�J�t��g�}�Q[�\��9��+;.$֧�ź ��A}���c���|T�xW�t0�s�r���{xrJcRD�5*W��V���oQ*�{�u�|���Z���[����Sw!���������G&MËg@��^&�"y���-�a*����[�9�l���-���a�3�rYC�/r4%��,2F�{9�����^��A��]��k|���B���HCM�2g����N��,&r�	W�,�=�um�T��*���k�uڿ�H21+[b����2w�yJH,�,��'Nv� \��ǖ�<J�#�x���G���Ȉ�6��yS�b�NZjk�4�`<���֡\|���yҫ��L!���7�l=�t� 'h=}h�V���)������{��Vi�r"�F�q����1��D�.���t[��s�N��0&
�\)kJ;:r |j�1CG�;��ݩDpr���f�.8)�3N�M��s�I�s��"�^���g�.���h��⸲۠�yo�{�3Jאm���9���ļh`��0x�W!�齎ܽ�dG�T)�0+�&m8�d��1
�=<^��o�R{1�������7s2������IfzؔS,�+*�?#0�L���[�[6�

�U��&Vи�E�'��im&r,|��TP lߩn�Hڵk#���H9�NC4oV��G�<��C��.��֍\�CLŐ�WQ1S� R�`K���TU���A�C�de����h��D	��孡1���ApC��Ǆz֖�$�3}�8d;@��S����I�۹x���!/w�w�U5�hu�Ή��'Mw� �Ɏ8�!�;_B0\	���e����"�@79��xA_��O����d_M%U�*�A���W�ߪ�oQ��Xb�mu���qJ�B�CEq��j?"�i6���|�W�������̛��1�B�Po��Ľ)��� 1�=�,;j�g�R:�-6ֻ.ER�)��f�lr��A g�t�f���I�{1<��������O��`�f��#��S�փG�7� ���܋=���Ë�5�� ����@'�`�d�l咲;	A�[��V��:�/3Jrhz���s����5�vL��-g���:&LbbTbI� �V�ƘP+��Y��u�z�ҳ�N�I3�:�[+F�N�X���I�Q]у��99�؄���9�(U!qm�S��R��^(�Y �"=s4Ȕ�#,�y�w���kR̋ћ9RN!�X�n՛�h#�IY�bٟW.h.}O��{]k;��!Ȫ�ȅ�)ި��c0��o�P6�.�,�]"��Z>Ԋ�(�v��]��	��Vِ Z�=r�sՅ��q����C��M��*�̔�/�'��X�?E#�>��)l�-E1P�ر��M܈�PE�K��d�|�'k�'����+\>9fC6i^i�W���Z����ofJ�Ay�C":�0`ؙ��`
i�$���;���-�βW` q�4����(�U�}�5�!<:�Z��K�<�O=
h���]��i�!+l>@�W �sI�dPmS��zgԏ�c�}!��'|f�2jLs;�o�����Z��|���ϼ�_F���l����;\��"S�����D�) w���fb�	Z`jLȭ��
�;��Sxiҏf��¹d���%�(8����z��{�"�����G�mDڟ���3� �G��]N��w���OVZ��e�����F�u��}��
�Lc��>�8�fm�@H��{��M���On7�
�ԏT�;s�"�9����]��J]�A7EhO�N��0L!G�mV�wg^�OG�I��:]pc�҇����FT��/+�1��vN��,��}�ϐ3�m����T� R��(�>�e��B�n*�wh�S��W�k�����v�I��ۈ�� ���"]�������e�����>UNþ���@�����>���9;M���X��O["�W��KMTG�J���sǊ?qH�?�xJ�~S��]B�V�%:���r���@Uȥ:��6��?5*��-։�$2����EG��%[N�*�A�KAu�Ҩ��{,5���Ta�)� :���~t�68���o�ٕc3��9{~&�P�qH�.]JL��ՂXGrE]��$UG����J$Guΐ����)�奲p�mK�d�U>c�rպ,N����� ��K{XZ�Yx'�r��6G_�J�)��?u��B��Μm�>p���F�]s5L���%�V������~�ȩ��n4��/�Ț�$7�!7�e"��L^Y0y_���Rd�������a�m��%Jg�Up��V۫��as�j�b^�1A#<�d�l��/D�������S~pT�x�U��^����zYj^���.lĒ��e[<T�k��6�
6m8�h|���YFi(�R�zn�h�&��GA��W~}	��g�i��k䚡%�#��5�� $��E�/��4�����w��G419����酽zW���}�lzb�Ye�F��Դ�I���9sgyᐱ��.������i+�L=�t�)�)v��v�{��4L����88>NWov�"T���(\{��9�O�]��pq��=�t�j_lC��{�a�}Q��
�|�
�t�39�U"�%��B*WG�̈�5��;w��@E�����7�e1���~�
�#�nN�˖�Bg�%t��F�P���] �5����F6vSx�~ ��7
��q�~F���'�?)��x˼+/h�Lx�a�|�~R��������QyMţ<2�k�`,^L����\��yu��������޶E�"^�UTO�"��Y9�ۙ���T�U��1b�$��H�vč���M>,� -&���FI]��]�j ̫l�-�_�{�d�Pes��W|L��������b�G�s{l]]������MS~~�}�.hMU��|�����/�s��!E�:�P�jۜR�� ���i� S�/E��@Dp�o�sk���<H���û�򻑜�ziX�K;R��%Q6���\�Q�@�e���m�4x��!q�[SW��?������x�}N 3,���أY�NǞ0�h�À�3�}�Ʉ{{[C���އ�Gv��Ѡ��@c�u�Te�و��%c��o����[j�Ss��� R�^7e�dL2r��/j�T�o�M���f(��������Uj?�\�����^c~���:�����ͤ�a��B0��x>4��$���MТ��J]��v�CN����W��z~��Gm9ְ�]B�g̰Jj���A�;؋{��T�>I�5�G��p��K�9�;ѷV�w���o̉	�_4�EJ�ҫ�Bc9n���3.t����7��P	_�6֯��z� ���	#Ef1/U(�^0���A/!Y�``�>6�=�,��	?�J�_��<W׶/⒛6���\i6K,�+S9����۸+�W����9%+}S[�!��`�cl�'�CQy�c���]��m�n�v��<\ �&��Ea�|�.�ĖE��ű212�1MD������{���'��4H�qa����aVRq�II	x^��bgI�����U�>��ے�S%3$����?9�X�펋am;����I�1������G�� ��/�Au�T��<W�7r!�2һ�n_;��~[�yR5R?��VÔ�B;T;����JtuK�O���L���aЬGE��F���2��`�%f�ٹ�]�v��ҭ�:�`��ɣLW��|�w��v�-fp9O&j#T̮�e8�-O�!��'�2��Rf-��&�1X,*܀݊��.�wl�q�U�¼7cT�9x�`ڙf��S���k{,���k���p韦c�Si������j��?�{��_E�c��5ُM���Yb����ڮ{ƖK%��n�%�߱�iu�MRF�wj���0����n�s��?ѢJ�����^����r�:����P]ܡ=Xl�0�Re%r��@��^Zb � %+l��ѷGY�ˍp�e�9w��sA�R�'~g����^cH\���½4��E_�(l���;�Ю�l3��pB��m�Ya�OX� �����K�d��(3n�;>��f\o|�J���6�z��-�����$td�öli�Yt�~�UC.>�Ҧ����cg�k�8����CL�g.k��)~F�eMG]�Y�u�n��F0]�F��)���1Ql3��J����[�|��dl��l3и7=��ɪ5�ݶ�^���V�ͨ� ���NH��B����w?�mue� �	��IU���ݩ]��n�T;�f��i���Ʊ�3�2�.{7����BY��k��䓸�)����u�K��q�/�9�_�k�
3T�>sJ ��F`�ր�Ue��.7�C46�+bQb�+-����ze ,�	��0��)'���t~�8<2NK}M��p�a���6a��.7�,ƅ��m�����?�%�K��'���u����)<�Mx�R���\�U� �G��!�u�8���%�d�[Ϣ��0ő{H�2:q�����`�L?�WCi��N!��}ZY��Lț#�&��M
���'��i��;�����l���{Y��R:�7��U&e������G���b�Ɋ$J񦷺��\�Iٿ������/�~d8&5R/lR���q��h�|�6�k ��3��yT���+m���/�44�Z���B�*��e�	�t��N��8Ň��NJ ��BN�H�'�U��/�Lh�.��f�rt.�\2�1)�:��Y#�%P���
6G�.���N���* �b���2���/�*O�l���e���	<��Z�9�ۨ��l�aw��c>3������L��
��^ҮՑ�g�ʽ���i1�=�.M����K/r�;2G��[O|��M��*��%�z�¡�X�dS��
�� e)sY��V��T��6�`���&K�flZ����%_��d��L"�t��瓕�)E���&� ��z���Xi��71���r댧l\3sZ��)�tJ�Ѐ��+3�����ق�����]�zlrHw��ۮ���DS-!v:�������n�C���)~���?:pǋ�p��f8�����UN��@������������@yRK@i{)����c�D/��ؙDôc6Kѵ��\õH�P캀2�����'pzT�� �7`�����8�~BƔS#Q�Q>:���Jl;H��)5G��D��װ������Ҡ�h,��,�Tտ����R>����+{V�c�K4��V��(�����P2;�To�镾��A<7�;v�5���8�w$��R[��s��1�gW?�(AL�Yk����ɶE��Z����U�"FK`�f�]Ua}M��'�R�Gw��W)6t��wȵ�G�g�a�t��f�.�R���B������F��US1!J���{��l|�VV���0�������)�t�&vu��k	-��� �#����<���g�JV����6��S8�2�h�b�������,H��tB��o�'m��E|{���������'$�q�o�{z�O-"�����Uc,�"��
#�6��鹞NL��~�z-�����غ{�eTP���x�ջb�Zn�d�'nB*Wɇi���ˊ:�E�*1؍M��1�A6y�����#Rw�� (�`WwB�J~�`��f�
���3��3ᾎ9������$�e��|A�[�jdV �op9�>hE���ݘ���dIi�-y�?r�nU���A�o�d����ZohT�����^����i�@�2�CJj�4`��8r��Uj�V�#cT�����/s�RcT�Hˎi�r��=��//����Kѷ�7���?����׀M�ާ�����1�R�loz����|xO� G!�3}Qͷ�@ۼ�Z���W�ؐ�������Sѷ4�˛�U���{��e j������] &��_��ޣc�'�u�Mw����+JJ��c��3�~����-E���YO�#7�4�t�9{#\���3p�_c�0밍l�Lk	�<�;:�T���+����^o��"]�sÅ�趥���%k�Q��d<�9�l�h���z��{2�{�^3M���B��0�mTrL(�S�GJk����(@Q��42ط�C�*��d��H)�N6��<Ac��!л��_^�ĺ�V3�}��I�Ns��,,bt�5�l��E���/%P���6�f�h���ª�:y����{!��7�|�L4�eb�5�R�MA��up{/�¬����ɷ�0�K��$�bYҷ_&or�KB��K���5��6/I��Q�{��
����~�� ���((�����(,[�����`�+�4��"x��"B�����8Ť�~��\��f�;~���̳WQ�;ܭ��7�Q4��Em���j]�eW茡�Q�S����-͖&θ�aҼ�2��Q�i�����gy��ū�����:�4�L�F��v?�Dp
UD��v席�+F
{��f�5ME��$����8��g]�'U�P }�j�l�x/��)������1	4�/��RN'>_.laP���%�>ҋW�#�ǉc�x�%�0�-��=�E�!<�(@���]E�8o���|H.�`t�T�c�PiN��b��X����t0���i�[�"1�1�9�7c�S�bl�`fN�⏨�N���ܾbD��t��f�C.���<��L�UC' 1��K�ox�N,Wfx�B�p��v^z"-���V��x�ӷ��-��h�B�)����+�g%I��Vj�7m���%tU��U��KR�S�+-&�%b����T�ٸ���	��Ã�f󞲂9��	=��հ�%s��r@jg�����z����Q�Wp1�������C[�A�7g�m	�e�tź��S�R���\x����-�yB 	��"/�iU.���]���~h-CnĒ�ً�_ŒY?I9Q0Y��GMASwC�fyl���fA*��K���wi)ɐ��d>��I�Ѥ��Y&�����<�.B�z�4��q]V{�A��@x���)��q�tQ��a3D�F��`<:�j��h�r-~�J�W�h
/�/��M�~>O�Ǹ��r�1a�<��b�X܄D�:�"A�l;�+Τ����S��:\��Hg.ǫ����AFH��my��η�uK�V�2��T�����Z���L�W��Oh�K10����) �
?�H�#:���\�?sFQ]g����&m�V��x˭É�v�u�Ĵc�2���Yȹ:N� ��A�	��P#��n^k�(����,������)��J`җ�d9���[�_��Eٝ�}m�y�v��s�8�ץR|�9LC;|g|��g'����M5�@�һ$�N9}>p"rD���XͰF�l�_o��f���|���-����[���9�.YWK\���Ux#%�>߆9���8ML�ӏ�k{]p�PE���͙�.���I�v�P��zs qe��%�"�SM^�Z$��lhc�Y�y(e��x�uD/�@�{�#�:9E%X�)D��P��*Le�
V_�������ۃ���h�mO�����WUbaZZ-��89��'�b���`j\^_���qZ2������f�Wd�EǍ6���(~�ii)Q�����y��ݣ��Jhd�ݞ5 ���G�~�0���.2�U���2���Y��sEv�&M�.
��ȿ�sb��"h�z��T��\ǅ�N���E1���C����j-vC���*���>�G8]��|ɜ�1�� �&	��#�9"�<����JK��2��C�$��4Z�U��.��Z�2:_���r�6#�^\���V�~.�O҆i��h:-u�0oEuDī�kb2�FW��Š%��l���ao������(�>zP��m2!�@��#���Fk	�T�M�V]��ȷ�����$��(H|0�/�Q��̿�
VcMW�_���	�t����f�����>��
����Jq$d��c�ݎE	z@��oG�o_V��-P�m*�6K�h���Z����λ1������6�̾��S{�����D��a#�_�ʘ�;7*������?l�������'4I�O}Y �m�v{�(��a����*�D(�B�P��,�G"\��<u�\�kѺ�yP@���|[$�u<�[0�v%��"jL#����EXϳk�b_O��.	ڎ4A[+Tx�)��ʈ�����N�K2vD:� -V�5�=��4��2`^�ނR8��$
�>\ 'B|�G��ɍ���9��#���z亭:��R��N6�����|b~���6�`Nk����m�Ga��qv� �?��5���}�˷T6[��JooU<E��D����5G���|�A����h�x�Z��0�>E$�7&�BL���
�Bv�6E��T���y�>酚�W����"��0�fl>�<s��*���sG�q�en��I�r�$��l]�l�w�����Ͱ��ެ�5~[q�hY�J+��y�w�1qfu~�Ø��%�ZDt6�! ����T1�����F�s��FGUe�jBA`���Ft4#g���=`�p醑-S�,�r�ٱL?)���.�VQƼ��M��Uj�.���S� X�&�����[I��Ѿǜ�'=�H� }u�(�,��v7�x�r�F/��u�:��/?�1����0���|>%βX�d{��6_�{��r+-����Cu��:���X*��,��9d�<6fyQEU �6H2�\"IfE��J}zE��y:$]�j�ZAl��a�~�L=�Z�z��M�jvG��nN�A��@D����G��M�l0�QJ|�*@�h�W�� ~hғDBf;&��D��b��˫���E1S,�GG$>01�T4���^�8���휽�U��Μ�Ty=�8���
{����L�/s�#/��n�$VS	8fF�\b�c�N.��0"�W7i'�1�_z,��H&��Dd���3�A�'�G?P���1�xo���@��#������|G��恣�0��Ƭtc)\�Y �Д�6�l�}�n���4P�LY�K�a��;�]�h]���	�3-J1cL�D/ȏD���{^\<�k��:�Hӑ+�Ƹж<|7yjB&і���1���8�L|x�nbu��"����NT��΀C8�8�k���o��tB.�*���Ұ)�sh�����qx�����@>; ���p�¼QvdCh�.�ˈ��M�����`�e�|��s(pt�2R�S��2<�����s��;�����h��� ��W�ZUzM|�c��nx��Ju:��8 n]�T�(nhRZ��x�dN��L�W�@;�l�6�GEn.��ZQ��$�}͜�L4���b5"�AkS�=�<C����Ƌ� [�,���=�_޸[Wܬo'����_z�qck�
���a-�w����]Q�N�0����0�Y���w�YN}���uGR[^�G|�!���|�2��gX���b����F�yTgx=��aezrl��d�(����%��B<��٢%p��8�h�a�"iR�c��F`V�����V��<�� k�djDS��n��e��R�*���p|��9MX����);�(
)�{j� �&�|��5pBTpP��׏T#0�E~�.._��0ae��Q\]�o�`A�z����E;�Rq6�fˆ3�BB���vǆ+Q�p��$��XK�pa��S��X9��{�ʄjR��s��q�	Ll�P��PM�9FU3����1(��[�:���4�����QG�]\_�����5��߳q�!	90��4����7�Ϩ�Y	t4uL�e�4!\�p	�z���O�k�|�3o���zA�֜� ��/	�.������/AF� �R)�:-i��w�`� 3J�bu$�&��~��nc�1�"�eJ\.ph`RRw]'��A���׏��k~��1V�Ke�G�[
�����>��F(�[M'��=C��(���5�I'0@��.p��S�d��cFj��c�/텕�|m|F�m[S�?�������Tl�ۭ	��o*���_<Q�b�����(IP"N_gh����I+/a}NC�6f�� �jvg\F�m����	lZ�F*qt,k�'�sϠ�a�b�s<L����z��w�B#wn�<m'k7\&�^
gᡴn,�����<Q����gF�z���&�����a��k�BIf�����@�iq���z/� �0����1*�XО4�\R���-�i�j ��U�&r��#����R*w�Y?�E�m؀���hldF�{��c~�B(!)DD����
&�1'��ѹ������?�U~�ǰC�S�}���!��F�����ܱ7��#iQR��h%�DF�cop!x�����M��@@��	��k��&�������D�A��+}ҡ5SS����	ʘ���_�C�~\�rT��c�M�K�R�~����P3����by-���4�Fwy��Ȇ����&�YZR*5JSG��x��i'a��W��E�s��W���	r'
�&�g��b��[ġ��l��Rd{�rU�"��m__���-�5L�x�����((���_����Jn�VV�YH�=/b�J���ǐk��z,/|ׇ���������A���
L�j��#���P�-g�o/���*��.g�G�J&���/�0�@��pH��U�<asՑ�]I��t4��a-M�c)1B*�y���O""&�`�̳F��iZM㨅�#����G�JA�|��yȐ�ޠ��=�~�x�d*v���L�2���V��'��Q�L�X����&��Vۜ���`�_k����a�wU�X験�R��B���y!�^m�B�dL��؜�T�6~����B9hj�	�u��bf��{�	��VO��6��\w�^v����bQ}�+-4��v�������o�j��ۧ�j򨟨��� �����H���R��d|1`Pw6��2Zޱ�ڙ0��?�''�Ԓ�y�����o�����һIS���I+���'�=��t#��^�rI��r����|x1���:ˁ����:�m�Qp�*%ZDQ�����v�!8�wu�TG�h�^�@(Vc�L���r��Ђ��8�h����RǌS���0����O��+s��i�ukt�0�d�l^"d��>���#�	��p!<)%A�����'~�k�����̡P�����C��Զ��$b$>� 92����^���X����o���i��W��l�_l��#gD��Ȳ�ΛWt�P���>|��Π~��XMzQƾq��>�w�l��8��Q9�`��R�RM�\�CZ�/P�ʖ\����e=aFfb��qb��d�$��:D�L�==��ppGY�9]��23�(��LS�ظ�bg��UHĈŀPWy��J���k~۶�huB�g�*g��@.�]5X�q� ��q}��m�ո�v�Իf���CԅG��m�WR���H�Т<Qd�� �g�nw��$(j����f �'�-a-�$���t�O����%�Q�n�@�X��,tZ��-9 z�m@�R���hO8��݄vt4Ɏ=F�4���;Ds�k�a�1�R�|�μk�z����P��B̍��4�����w���4�+Y��T�@1Wz�o�t�^ڴ��b��6�fص�~%��lD�qACQY
]��D��L/�ʳ{��!�"E�����[ϥ��������l.�n^"�=k�@@�3�~=���H*�-č�c��ԅCz��bAu�����gq'��i��Kp%2�6��+H}�s����d3m��%|�J��i���H�[�Vt6��To� ��^�{��,A 4v�����J|��L0��&���*p��yf��x����6m+3����u~h�"Z�=eDy�{��R���"£N\�l��B2DN�Ⱦ$��}>fi�4g���MNF�v�rV������t����E����{� �d��,�sm���d�D��eU���%�R5$��z<[�Q>o-�̿��Ez��*�5E,�G���:�����`7�
�x�k�nw��v���@ j��B��u�!,�O���w�@��^��P���J1��;���4�����aGP(����M`���ɍR*;ӛ���8��%����Q��m�8I�v� ��ާ����γ�u0Y����-R��xS�xx2ǽ�T_EC3��+�>�
���âTp%T�we�E��(�(q�~\������n�
�q!���W�49	�p�mb��%ޜ/�5T�i]&�kX�#������pr����sAp���*�ȹX�����D��'T(��N��lJ!�ǙhG���34zÂ�i�W+4��Y�E���:�H���m���|~V�;��u��g�]��H00t`��[l��n�v���̝���Hu��]FlG?����Ю���#�Lb03����G�\$�uS�n�8��#%P\vs�s����E��5\0��]���?EP��� �����2�P��g���O���ěǩ� F�n�x%�ǎ���O�!�d5�a�p���t��B�qCp�@ARaʣ�G�{B@$I�r�a�Zų��%*xɽ���ٷ/�-�5�8-d�޹���X�2�N�[aw�7�1oKF�(�v�R�}�z6��T�TI
L5Td�Q�Wq��������rϢa��5��0܈lw��$Da��ѲP�B������Bwa�5m�H�J��C�t��
�v��m��uN�����Ӣ���u:���}�=�)9����66ƾ>s����FSx�r_�q�,t�%_ %+/�3a¼?X'5e��A&���t��%O�L6����%ZK�z����*���NO�9���m��J@�¾��`鬏q�/����R���l��	���Tc-f>�*��\��Ք\�Izx��T�����w�d�����q0 ����_:a*G�Ł D��b�G����0���Ƅ���IP8xcx�lƋ}��HH��%w�=G(n�.��c@[i�hG�@�	9oA��A
��=ϳ�/���8�\K�D5�;��;�Չ+��i�zj�	�ߓ�Q�ax(�Ѹn��^Z{r���hW�7�\S�\��'픕�/��"�<�*��A��	5����Κp]�!�k�3��o���!�2N$�ٖ���2z�cA���6�	6��	���"�{�7;�r?����G��9Rg餎d|�mM�g=t�Q�(���/6w]b�t�(���%�&_�����U�ht+h���<$����ѣ� ��]t��'z��Q��-k	hB�����A ��*6�QvcM`Q"�&	��/tK��ŝ���{�wy9�nH�Sϓ���Xv��Z���V�Q�<s��4��s�e�~ɢl�@0�	z��P��qJ�6E�����a�Y�B#:hG��@���,���eB7N���<�oQ�m%�v-�'�:!�����ߪ�1C�ߢF��9�l��oS����]�M��v��I+������5�_����)�p�h�9 ����hn�c�÷| DъL]>	&�o$=�V�){��gC�8�f�AM[�h:�Z��A͂	��"����FpP$az=!6~�!�5 J)m���n�ښ�;m ƄП�]Q10�Z_FݕSc�y��M�#,8ȸ��ƶ���nn���@\�@6g���q���%�er��m�4����IBV��P�PTl��҅Հ�,-�չ}*%��^y֝ID`̀��C�`�a��y^��*���Ӗ"2w���h9O��fO5D�ʃn0⣖&�0�-���#��'���-�֔�����j��.��D���o���h�� bq�ޱ�t�����KA�L7l�4�"g�|JL����"KX�~@w��7�g�X��d�����
���A�ß�GL��+���G���RiP3�-NZ��������gcK�dɦ��V*��R�+3�oo�lqf�)�t[D��*w��SVz�W��o!��Ky��[��E	�z+�ԫ���kt�Y(MD�#M��)��s2R-��9u>N �_bY£�l��&�
Qx~��R��~\����إ�:�8Y� ��х� �1��j 0IH�����j]���(DuaW*Sxf���2��U�d<v��ϟM(�T�9��������v���E���
O�|Q�](�K3
�/�<~��(b]e��(?'�_�u6U�G�u={���ȳYj��Qr=l�\�2����D��@M�{6�����g[՝�2�JŅ�2E�2���0�+��.A���ꀡ?r��Xf��۫M#��k��p�e/�ȃ�@6�)ت&� ��I^T[9�ӳ�A)E�D�и��oR���ל0_^0^��#6�55WcN
��0F�(�"����K�ٺm��rM�k�T�Q._�|����Vq�3�����IK����x���A�S��,H_��bO�Е���`���<�a�	W��͸j����}M�Ϭ�J��kc�Z��#��ND��4D����"Rlu�J��N��%\�@���G,lf�d�9�Q�������t��7�m���s�z׭"��q�)�K�y�d�)C,G��P�����j@j����&!W����"j���zd�j#�i�[J&(��,ף&��*� 03MXe��4�9�����^�b[�{��`��ν���X��п�N���H���lf�@�w����Q'��oi�?%`|�h�C���� V�J�j��?g|ٻu��OM�[�֔Bu$_ԥ"k+��,K�$�0�z��t!W *狜�>J&x��!p�ҭV�5 d�_D�׭w��38?����q�V' ����+Eh"�,�� =]����b��{r�d�
cоK��,�T�4j����b8����?�˘[��*S�&]P�{E[-_|�&	�=�1e�1%�L@ȉɣ�%=z�`,,���Ѽ���y����.]�i��ڈwP���<!�`YM�&҂����[5�ʫ���b�$�-�h�M~��N�������0��#���\�w��K�ԏ�r�:���f��{?�p,+̕股���_�|�9gk�Te�s���"���/������g�|-%�+�g��~ƴ�+$�/����\����ș]�f���^�?l�v�vJ�F�����h���r$я��UUإU� �zY�Zӻ��^�K;�W-ZƟ49��_��7ժ�7�N�(������tY/�m��)�@��Hg`��'t��na{��솇=�	#��M��L��+�>��\|a�;�����זV&R�����/:Q֪������b��{���A�"-�y��05��I���T�#�A�T��&��tbH�o�������B����}�D�+�|*]�g>uR]s<����E]�t*��..g�'�z���B�"\�YUO}&;�Q�`�Ƹ%P+ �m�ܱ�Zފ�@A�+1@b}ʯaL#/e��--9��Q���4Aa�5�@y�:e(%�ŝ2���$�!ruB�}���&c�j^�n9\ȏ�M� Ҽ��we!�-���m���Byl?������%e���$7�|��'��|!����ʟ��pդ��KCM�i2w��(����� �q��~hT��~>��,�&30��N�p �h�c0j_�G�|Nek]0`����'ҡ���=�_��e��r�	A�x[:N]$ ��Y�q\�v�+�5r($�G�&���SMb��d9��*��N|/�\���ț���o��M�@v
7�r�|���N!�R�c��'�nY���Rt��l}~�S�0$�»�F��$y���@� .{�h�HO��4Lp���|Ȃ+����TPe�¹��y�g	~u+s�F�q���"Gw��}j\@��5����]����kEs
Ţ���8�4���I�?��� ��K�ն��E�@M?ʎ����y'!���Sl�?:ƵBOi���y6�s����S��z�J�P��?0I�)��������`��-t��jQ�i������L�ý���pv7׆�R<5e������;����A��K,oh�{���A��z^P�½ռ��bj�췱3��X�~�9��p�[En<b����r#� *�L�"t.f >�=��I0�6@�ϵ4�	B�	�m�W�ubࣩ��{�2�s=�%���c#
�fo�X�6�^�������x��E�XS<�K1"�c|�&�]\	;c���;[<�D���K�S2!�Ľ9��(Um踢a�mZ�(巆2i�ܢ~u�̇��+Up��~�"o-�����^��h��"z] &ݰ�F.��.(ĲDۯ5�!�T'u��4ʜ1q�n+���?R-N�����Ŭ/���6~��1
�Ժ�#)Q���a%�K�Qj 7l����������o-�R}����cl�ޙF��8����R u<�����==P�I�S[{�P��}j��mdr��b;�WQx|�s6���#]���D�MD��s#�GK8��ؙ��_�u�Kw(�h��0�J��l1J����[�Iv�)�0�T\yFP���G�p��:^!����.uE�����5�ffG�<��x"Q���)����f1�ĉx������6�}zȬW��{I�B�-H-q������ֽ&��}ӂ��Ŕľ4�R Sa��=JWc��9Թ�}�������0��qy�����u5јȽ��$�?5�M�?�(w��AJώS��9���
#s��k�#H�������,u�#��,ڽ��Ԃʋ·�dKc��:\��W��N1G#��Y5�T�@%�C����ג�vȢ~WD-�i�@���g���WQ�����G���|b8���6�EO��vX�wy��㣷��%d��,��j�^](S>�8`�F�P�1��k`�X�ۜ��!���|�p�M�ډBm���/�C"��~r��)i�R��:�\�/-5W�&��7M˲z��		����j����Iה@�m�jcQ}�mP���\ �UW�{�y�ԇU��b�^N9}(�`I����%r�y=t6X�e \��eaOTl�0�d���=E:d���\��3��VFfpX�}=�����|k�UQ�����o��2a����U,>��~�6i���b�;�=g
�P/��_����,�)U�P�{�.����au��X��)O�˕F�}n�^}ו��nr��=Ю�24~�g���:�r�N�w��xTC���H��m��/���G��&��&_h�ൺ w��[����+M�p�Ң�V���1~-\,�&F�Ϣ߸��z��S]��;��Űj�W�j���o��㞗k�,��,-3�3?pS{�=�ϧU���qpG�n-�א#}�Ib"�'wtU�q��w��m���
˔?鴢j� 8�0��h�Sـue���]�}�^�����1$����ݾ��	q���3��=ܘ<�4�d6SA�g�ܽ1�^
�?��wTZTh�o�P�F�X�)�C�k��,(ht��j��X؆�K��;YK�Cn�V|r��?!܂�(^".hH�p;�L�hmv���[�tRϴ2�@b�זX��Dn�SGZO���U �3.��_��b�Ps�k1S��t�.\� 0T�\y���@+x���ɧb����ڨ�y�LԌKB���
in�����b�����k��z�=�Cۍ�{ �:�뾉
C4@?�R�X�.�u������[㫖��8�(�)P,p�q}0V��L���u�f��&!]�a�������o/-��b���E�����\lƓ���ң�饏��7�@����&jW��5�A�%�V�=iP����֑�o��4�1
�W���8�l�:��כ������(��# H����c���=�˥	'�U��4&��!L�䭊1A�?�`�G�J3��o)��\E0H޵m���ыcO#l�x�G�V�ɧ���$�����hy�=�)���*��N{���̀gGj��{��d��Q��뺌�8"�z���2f�i��,8Cߴ%Hz�hvF܂"{UB�{<��A��{�����2�/���������x��{A��2Y2���g�e��u@�F}`(����q�N��u}������:�JWE.Yf��� 8鰦���6�B	I�[��W��A���[wr9PHX:��b��ێ7�yrBX�%*��9:`Z��1�����-�չ�+#��Cݱ9�_1���'7<PJ�'!2��6���fЌǃ�D�|�%ֿ^,C���[�]>��Sc"�E|*'�1U�	���n�V�{-0��[�1���Y�Z�%�Ex|�J�B�;HB��2���gp�[#���c����3�W#��9KcZҫ?�������/���ѽ��A�#���7�C���w����'Q���0��|���c*n���!��X[�B�&�_����U�����}y��|>;57�ݙYc}������P�C#w�e4����Ki�q)�Q��CS@�(Qw��,p�"v^�������nb���3�Y�#�Gl����7k�CR��W�Y[�1`<��Whß�W�͏�X-:J��3X~���A�S�uE�{����$�����Q��B5(3����˰�zEG��7��4,d�5Bj����6�KKf�E�Ő��� �O��5�G��>�~Ju劼��#�_.�}�`��P��Ҍ`���.����k�ݷ��ψj���9[����TV���0Uob�6�'�|~;@�q+x߹���.�|<�Ênl�s��� ^���eTgH�f��a�Hi����g*�Qr
���� 0�!���P��8���k�u[c;�������� x$**/k�"bN�U٪ xOT�c.F�W�B-�P��I2���^�kִ-�Q��))F~�۫�1Y�l^X�kd�j7U�T��&K�gV	]<�M���=s��c�y�^ZR��(̅�{7�$~Ϝ�G<�vy'u��] ���0�.�����0J��&�J�$�0�r�^�m�X_�ff�_'�ņ5�+)��w�|H� ��DR��8�)پ "�^?���Jvd��(_1�>���<�IǱe���zEzQ �~� ��֏L�q�~w#)b9V�+!�֞��D����Y2�_�>7��F��_�3?�Ʌ�I�S�8�ۛ:����׹��~x�ڽ(_�ɇ�3_�Z��'��ĉx�BŧD��K�CX��x-��-4bx�h�o]��a����$!:=G�P{��#x%�#oMyd��c��9����1_��*.�4��"�e?���]��� 
�f:5~M�Svw@���Ey���}�~��JT���Y���&�6��.���h��WЉ�V���!������$'��j)Z>�Q?>Yx�NJ[�j�?01�A�O������/~d*[��]�z/31���L����M1���SPzrj��ؿ����!x�m Gi�g�S�M������Ϯ�_�7�D�/�iտ=j��K���B|'3f3�H;X-�Q1 �r�w$��, *TI�����HjJ�QF��ZnM��]�D?G���:J�"K�Wk:�Л����H����TW��=�΅��������?G�	N��X괴������nh��1�q`Iv@����vH+��Q�uao7��O���ي�����o�t�v�Q�І`U�ω9Q&�E�n=eVU��K�P�%
�u0-�o���s?(�؅Н�̧H�k�G��ʵ.�@ PkGf tb��d*�g��G�V
���T}�X��v&01{�����EL=���k�Ե�=��0>��|M߅1�����"<u�|1b���f���-��>� �hpB]mRu���Z.���L�|?��Ⱦ�"XO{,�;G��Ggo�b�3�*櫪X�r�Q����!�;�M��Zq��B�5�Mc�q���Cju�_@��O�qCN����BeUz���x�+i _�$�Y��?zVf%��:?�Ke�4cpn��Mvz>�(f(ӏ��[j�^Քvٮ���R/"r�AgU`j����4e̅X����O,Q�0�� '�na
�gK	�/:8����
v�q�� N��Kh���C��]��uf����:_�¹(Ut$��$�?���3�v�G�."
�G;؟�k�#�{$���{ #��\�"����=C�` zS����0��[T���l��N4��v�u�������vު�fxl/������u� ��2�֥�{m~!�''s����� `�r�\�&�Jf<�r�t�&v�������6R! �V�[��l�+�Ӱ���4�"��� !�@v�l�%\��8p��ʤ㔘y��$��&�{�!��W��x%ZgK��f�Y��1V Z�M�N�����*t�L��\��3%���{��M/*̈��r�<,��jA����e"��h��L�
�~hU�듧�!��c~�ŦƋI�����t�	���s��q�B�-��}'�!��W�����W7�"�����2�����x�c��v�qH�����2��x	=�B��)A^_��RJ�7c�z��Go�n\Ŧ��<��"szј9�w3p�90�îA���e�ElcW5�R7�,KTC��Q��فlTxһ��?��`NM���
���^#�	Xi6Q��I�'���4�z����N|�i�S�����N�ɐ7�/Dc9r�go��j�%Y�+�~C{7xrFٔl6�E�����s��Z�����|"�`��.9(�F���gM��'ե����4+C`�!E�f����g�ٮW�$/�����
z�7���H�[��{*�{j���ݤ.��m�	��̖Sm	�B�����A���C�#�f11&���=�_�	/ڵV��?]�r�Tg
8H��-� @G>�\u�� M�n����:=�:Y�0�(�m�C��KǪ|���}�z�x��9�$�>�ߡS���(�aR:ݙ$4������N_\���[����%�KiB+[�>[�O�f/�m�q��5�G9v�k�Eɒ�i�ؾ�nC<S�P>[8�
��&J�WѱHX����3$���nTt�ƅ�&;���X�ٗ|0�h�Żvŏ^��k0eO��/D9�2���n]]��{��ђ���5�.P=�%���){���Q�����~#�j��:k4�G8i������2�+"X��;�{��v��!"/w��Q3um+����3�a%R �,���g�I6��Ŧ��#�� 1t���7�l��]���f@��;��L�Oѳ��T�/N1�a[�2=�Y����)6�hs��Ik}�vt`��󟝂�z}o��uR�g�v3 #Vn���\B��S.�`�'����(\�~Gݲ����WҞS5�eȅ�P"ʐ��'�疢�J�1�����Uz]e�O�K��ꔠ�1.Ĭ�ϼdA�]�ѱ�Q�B9�AY>�v2~.|�ge?�Iq�WSg4"ʨ_��S�V�zx.�� ���DΗ[��T�9���� ;9�>v{�Z��5F+�r$�R���OEﭱ�[�6~��B�c%�5=4�O�4@]��9U;���X����U㪢��Ly�fi��<����t �$z}����1����d@(>��7Q_����p3˛F)Q�o�|<:!A)繬nی�+�a�M�K�<'7 �=��tN�v�P��sȉq� ؏5�ί����b��}�@��p$��;e$|剖;�Wo�*f�M�e�2�n��@��Q��nD��x��u����8ߪT|�~{R��th�,^��x��VOʔ�pH�n|��8��P�n�!�@e�w�4���e-rr��4�`6!Dd�����ʪnBG��W���55���Qΐf�Eő���T�%�tk��Y̥���m�M����4���3ɤ��<Qv�_�ޯb{��s;���L�`�F�ͬU�}Iy�d���>bp������Jns����THߖ�H� Y���A�R:d]�j���3�q4C��`�S�Hi�
E�jrwpu�!�rѴXhʐ�Xaa6�6Z���l��=�.�[�~�e���¿y
���?�yI��ڣ��Q&�t)��ʐ�sE��&�˸4�=-��	B�Q���cz �c�L�8�@Պ�&�C}bn_ȟ8���X�{샮�t�M�R��Z�J�O�x�69'��1��݀����h���aX�Ҵ0�,��˅8���l�h�WA�<�3�I��		>n��,]��~��7Ď��K�If}+:�1&��s��<��
����\�Q<Ȑ��3�e��v��l�����ޙ���<滆4��B��/Lp��;C�0(.���KB�lo��@��8������H�*r�A��t��G>Bo�(�kv�E��_7��[������c8/�;�'^�����zSU͏��ۈYڒQb�퉗`(	,x'��.��b�Mc�OO����,�$�|��ɷ#���i|,��;FiU������L{�}�m�'��;�m ��/�7�y#���5u�U-T�1&��[tB��i�B?��S)�� q���U��u�bN*`f�P��-�n�~<�M�<��������$�5����CU?M�W�ٲ-��<|����?��<�-?��ȍޚ@|��yE��l�#ӏ�����pb�7��Kd�q�j�B�I��dm_���Ӈ�1o������D`�Fó��Vj׷���||�2f��L�X;,78�$&v� ]&�+~�n��VP��ꫢ�/?��2��Y��X�y��>�\0���W�M0��:h��y�G���^4��*���'�#���J�4���m�(���j6܋�duu���MGu1��A ��X�o�����"t��y�I�(�[���3E���ˑ,	u�uE_����&|�g�	#��c��p��4��1@��-\)� �f��g'�YYr�;?���4�8�9�B;��t�2�8�)�i��}��7��:�h�r:�dx�����i]�)����&m��?<����	Q`P}���#�]N���)6���"�a�[�+]Sb��B�P�svJ��q������*C�H�����AC�Йf�Ψ��n���QJKy%^aC����d޵si=ۅ�j{`�v�0�
�	�߰��F�+
+�.bh�s~�hC4�����-��f�d�a�^G+�����qcY�(Mb�?�J�J���Bb��<<W�f+[�>z^��.���k�b��o�ڨOe�VDI�K��og��� ��c!A�pB�U�s��.�����괴ƍ��be�ה����oc.`S[�K&J���&`�2Y��x������d�z��ƔТ\�Rr�6��2�om~'�H<c45�8o��kgj<vʯE-��c�M�Tz��e�CЩHT�Z'c4��[C�ޅ���vR�(����r�'�5r�ȧ�����u��<���R�"׀PVb�bj������t�\���޹�@g5���<�YY�%�`>���nc�/��M�e[��ۻK��)������L��k�BZ�O@8�nx�9�ڳh���gu���~�/��鮇l��e�V�Oy];�����%�_T뙉^t�q+=H~ �@C�nzm���x7]<��6p�F�(����E�L�� ��gO�Ϡ��;��0[&j4h���OꠗW�ɐ�T��⊽�LY.X��r��ܻ��}4�0��n��R���K����k$ԃ�P�دޙǂ�{����b|��Y?(I+F���J��2&�d�>G3<���7a��6�ώ�9v9D)�.��~|�Si뵭��6�GWW�1t�B3+�Lp�E�E'xĺM+��9�.�u?1�답f�5z쿥{���?(��o����� g��<]�#��p�P�7�;�7	��4�NZ���ot�:��$	CD���'��`Z`�����&V5�i{p����D�-Ѓ��*>�F�z�f�	���1��>S��E�x�.��ĲZ�Zk�tbВ$Ԭ��12yg7T��z Ṕ9]�N��"����ZF=UU�/4��� 3U^��m�����a!��|��&�ƲJ�J���D���1桱�<p������bX���S�p4�P��t����r����S����K6�du�v��p�x��B(`�W��;4}�)]�lAL���K��G bc���K@D�L9�y7���b�v�"�ֹ�VBZ�x��%���wmx�]�W�T0��M4�k�}�������ˮ����_�#�7�q��sV\��ϼ�9HT�zI8\���ІW���A�9|��}M�T~!�ק��ಹ:���}ʲ@� %��H��t�k㠪�8�����Oi�Zvs��	����N���"b�JͲW�X�����*�@�0=l�Wfv"��>���É��y�b�=
��������1 �Kg~�MW�����o؄<��d�{}룣�BU[�۽�qS
H�S�Q�m#��d���e��PSġmOj)@茸��7�S�np̒���o'��-�ɤV�|5���F/��);�����\����Q�FDz��5>6��6�is�� �_��D1��~�,��j+o��j~��23��"���
Y�ՈP��֚c���|u
tdgrK��.M,��)���=T�J�a�S�{z���}�6,����&>�~��<oq��?�۴����%A��S���Lj� ���}��wK��Q�Ȗ�Ⱦ��ep��+d��_3����u� ,o�����t�6�#P��P>��P����֜[ߛ���	v�2�M�Є)Du�I����\�Lo��%�rhh �`8���n6|�" k�5��:��iC�I���hc9=�C�1cQ� P��� U�T��ҏ���kB��ӻ-� T1���1aJMO������[eU'L$E͵y8�i���#��?lꇰib��-FW��ߤ�1��&��g헷�6HN�A�|��<IAG�'��D|&FyK����]¸ш��c�߱�-���&+�+lh��SB�Ĝy�]�)tC[�<�	���?����I�~�j30�i��үc�m>A���o��"���w���PP��o��GE�\��I��3d�ݔ��D�s�ȵ���h\_�mT��- )�@��˿}Z?u��RY%��Ņ�U���+4�M7�,�a���|���}�71��KOF�2BŤ`�	�7#�;[�?:E�̍N��Z�(�s.+X�DGfC�m�N��X�[=I�H���^�r�&�6ef!U�Togus�ty6�`P�Ԫ��QRՆ��Iq���=��2p]��ؓ���<�V��_�A+Yޡ0���\���?�+/O��Tv�?�O�v��Ɇ�לu
d��=���&�x�Ӝ=�\��R$��������0��rw����� L�F��S���Q�)un�x��O��C>T�Ȥw��O�%\��C�1����X=�7V��������)?�^�h�E��~�&V��Z@U' �,{���ۆ\���=0ՙ�>�rx{1�΢�h0��\O�:����x����$,>`��'�9*�3�������g�ؑD@9��$��d���N}P���Y5��p�U=IQB�.t���_TW��'f|��*n�{GO�0�u���y�V���Ƴls�����d�>��n|�S��5<�|��Qg��ff���#��c���-R4Զ�7��`����ܫ�4�("��]�����\[Yԟ/w�׵����h0��ԈCd�H��3����oG;т��}du����P#?��KsJ��4�
Y30<����h�ZM�`�[��A��hKS��f����7������[�.�VL�AqRz�-��o;�a�ъ���UZlD�!�=���C�o�6���^�t���+��0η�W�x��^�vh��X}��e&?}������a�����rLi�.ZБ����^�{���:���k+��1�䂋f,N��Y�-q���	Vo؆|q'����b��4#�+݆ ^fJ�i��WE���;B��^����bW}� �?jm�h�<�a<��=��J�&a���k3��Oi���y��"���:���p��	{�D�/Um�i/}	9 ^[E�WF&p��>��;����wO���ܼ�>>Ϳ^�y����:�m����1���#/���~x"��f�&{mI��	��Z�$ޔ�wpGf���N�*s(��<�6����܁�a	��j�Nk'*� X���v)�-�߳b�7��F��w����S�y<=M�G��|��7������uFG9�|9u�Ռ(�d�L���34rE�%/���T� UΖ�q�%��Q�C⩮8��[a�ǳB�YP����֘C�x�"� ��l��#�����.��b�I�-��"���%�3s�� ���@D����>�����}y��\k�3���Y̗U^��s�p�e�vN�i:�ٳ�y��T
�$�Ы���A��ą��J[��;�Ko:Gl�R���d,T�h:���<c�24tG�'�q�i���ف9�xX&$��[��%@ߕL=�b�f�c�
s��e?�rٱ�F�v�z����ِP������z*�����/�g�5d,}�N�=����R\�x��j��{M�>��#�D�6	��j�$v�B}\��W�.[��Yi�!Ko��XD�v%Ud}��b�`E{.�W��9�21p��V���Q/�k��+��2�4��v�<����>�W�(���M����h\�w��j0�Z���n�WɥZ��)�j�ٖ�mM�3����.W=Hع�/��Dȴ�4U4���>��g$�D�Kx�iP��=4��:o���cZ_��I�E��\7�
��G�F��)E�Ei�F��n�m���
���� �I��m�;���WČ� �P��7����$���xo�C����\�B;/��#IyD�$���c�U�f�(���=|�C�iU���K	�V8>���Ծ-?����k��?J��.��mO�C���H�"���l3rT\��p�M��`�o$%F��<O�W�����%�C �/ZO'In:v��h��9�+�jc�i÷q��*��t����0CD�Q%QJ�a�;�L�'��CG�%��b������7�R�E�@�f�dB����f��j�z��ω�.JD���/���r'.��P��s��5!�kG��?��^!�g7F\��������]DPԆ���O}[;�O�f���AgBiC��0�%L��b�:��
y�i�s�`�ES���ӟ��%=��:-��?Z��^t��ܾ+��D{���]*��O���������A�n4�bϋ�8i�9�N�å��S\�-C}+�O݁�\M���@����'	�v�w�hf^,识��wj���]J����i[K8||�P� K�e`��r79��"�T��Y�CM5ccZ�P��u����)`��� m����r�әg�s�+��Ԭ:]2���B�b@	��Fޱ��g���Pr���0�j/�s_l �����e��'�|��!�{%o;�r�ID�4n���G)�G�g-@!�"�P�zǪ�0��3CTܮ.U����w�w�3c,��pȝ1jdI��5o���´H�q���2�+��&��B�]Ϭq8��1�r3fh�&]�*�pvfUZ�_��sA��z�\�|;�դKI��A�qR)�g�xv"�L���Mɤ��S������(l»K��C8��Y�O��of�����Mms`	�|���b�I��?j��(b�7f�*k̐�e�T�� �GR<;�=������U��M�[2j�]+���[=��"��ɻ��&��pO��˿�D�-�9[Q�j���E:/`;��2X.i�1F���ǥ�Mx���ܮ�� �� �� �v����w�����@��Fj�6�m=*�S!�1������/��(I~6����.C����;��&���{���!�a�ht,t�Bǲk�����oT�h�L{y��o��w~u���[4�k��_*$��B.Q׏����"�A��Y�/'"x7G�����"h�iv�_��D��>���R�7�gaƹ�H��W9�g�����4BP &K�����?Uޑ�ԃf`\-�t����C!)k���TH���w�.�`�ћ@w_�( �T��,_,�cϚ6m��M]�[���{'�eU�� "��W���`�Tʑ�y�"�K֦!��Z�q����	��E��G��
�����,2_������e�zj =;M�5b�FR̢;�Á:�]k����	*\���G���(��+i�V�ĽظPj��p�; �+�x[����N-��K=L��P�2 �!0I"ߓ��߷�������Q�*�yX��WpY�Ң=�,�ԥ�ܹN�"yF� �Br���*JN���@g��붹����ĘN�5,�3_�" �.UN�;_��Lqgc��i��C����`�C�/�j�* �5)��� >�>�5q#	`��|	���U��WcBR��%�*�ȴA�����P5LW�&��y<�"��<�wNt�o�9��;��<�q����.o��ȯj��h;J�z�~a��8�_�D*ԏ�&�[�0�w�0�\���AN��R���O�8]��ɂ��b��t�`�!l���=f�cH������e�s��l�k�6�����몌�ҵ�����;gP�`���'��%�2a��|�;p��L��6����\2���Y�� ��T�����͠D[T�J�g�ш�=2+c7x�\~c���k1�5iJ�Gc1S�Z�C��r�ʟ5Y�ͩ��o�#��fpӀ�M*ډ�'u9˂:rһ�SX~#&k������7u�׶�5�I�=�4�(��e8���7zzI�k��C����$ud&�,���{�"��g�)��MWs��Ջ�вH��v���`$�j�?^Û���6�j��=`o��ϒ��9tr^�,=��K鸢M���'����������xh>�p|#�e�L����'њ��69��<��6ۂ=���N�����z��,���)^��EO�]/����R��~n�ΪV�ANì���kϝ^�J}�L�;��@�A���z�9${�4�"�<7ى�]n�4�Fr�4 1�	4v��V��][��$�.�V�Rp� ��
�\�J���YR��6L���8�P�d��A��r�S�Q%Z[��8K���:�i'x���+��m2������3�E4&��b��2ǌ�n�q���d5����b-���
�>�kf�tb�J>���9ɜ\J��KU��'�7��F��7�կ����IRi�#��N�+����%�Ԍ:S+>���u�^Z8r�o�2AmX��Ďh�&xp>���.��NO����z�P(ډDp&�ˏk5ς���P������UFX��S3d��Bo��f*mځ����"ŠVu�p������ �s0jxY6T�.A8/!Y��VoԤ)ۑ怋����(�@�jO%�a�y_�_�*H����f5��/���&�S��WL�&�#\t�c��V�֩��{�ŢF�ge��+�t�����d-7K]t��ľ<��w�n�=�w��.5�u���z�=XO���pjWc,�(�i�j��?�X��J\��k>�j]�:�s�l� ��3�m�+I5��1��uǇȞ�4n�J���Q��cJn���}�8sZAaY�3&"܆{���_
!�
s�����g�wM,����@�y��5a���J�[?,X{ ̈́�9�����2�U�{� �����2��Y�/��C�IL<L����&�?�L`�|T���+��J�;�ږ�_�qG��2$o$�H���=���Y�mW��R�iKT˳w^�JC���v���!wo�d33�T��zXO�`{���'�i��0��
	�0��L�>2|2s���q����5l��Ű!�{m&��wj$�n���x��u���TEjO�����r��jm�[գ�R�lnF�X��̥6�!vO� V��=5�� ��Q1~�ݕ�p�\��58YJCb�E�"��V|6�}>a�dI+�?x�2Wʪ�@\q����GX	$�ת4�$���nf�A��v�?���Λb�K�Pr����QS�1��0?�;
�+��(�d���N������/��
�kȏG�װ���'����!����-}�����Jԫw܉�N.�ҙH�J6|��-�� KB��Z���� �=��&z�><�j��D��U���P�0�;��(��K�����k��z@w�X 6dW��	�j�0� q�Lw�9'��o�rW�^�qJ$��<�HlUR��e���#�>ḽ4-�0��pr둈�A�)�X"%�7��lPx8J+�EҢ���{�XC!�Lz��q��9�Ww��H4�p�^d��zF�Eg'����ra>|�����ɽ�Y^I`��T4oy�`��O{����p*K�P�����Ş���N�$FcO>����r��<�,��D+n
���!5�c�j,�[V��v�UP�.���+
���t�H�{r��=�$�{ ���n�XJ�H��mK#�L{Q���*����1�o��,�-]Jy.�'06H��c�j��V��3�ͥ��166�%�j܌��������W�z�Ր����I�'U�#5�bHQ_��)|�8��q`| ��kZ�0�jz>M�P��ձH�q*��E�o�O�<�`�B2yy(�G4=�&x_|�/쫕�S��r�$#/r����i����֙ٿm+������#{=�: $a��a�z�#造����^�#�8z���- 1���|�)��u�>�m�J�E4u�홽�H�p&�ak	I,~��ʞ�"Y:��d�P����U�S#80�j������<ִ�|�=5ie�'�tR�U�9���!����z���G�ύ5QbV�᤯f�~Q��82{�nĂo.Ϡ]���*��E�f�֠(�CK()�y9t���Ճ�S���<l|z�e� y7xA�b#��Ʊ�?U��vJ�������wjS몽d�މf�J�=���ꨝ��� a���*�����چsǘ����OPK��P��هj���@t>���y��:�ᙅ��P��w��qbmI���z߬'���_�ʗj1�p_m�nj�������h����wp��u���/],4�ɶ�f������z�yq(_@�X����"ڼ/;,�i�z���9P��'��4l�����%�� �ec�ۯ淋����4�>w�C_�n��?\y�S5��e�Z�7(����V�>jU����"����ȍ
_�uΜ��F�
�>�8<��B��1Qg��<��U�,D�U���n���̗���:�'���g��g��s�r�8���(%�"�?�����_j�=�O�֤O���_��,<M���	��~p�8�F��m�*�8�;�Ƽj��>:-5Ud����AB��J�+9��IyC��(�`=�UO��ᩐ��tˤ܆j�Ty��:�Gۦ�a�\�ők��=���s�a�ɗr}�Dݻ�����n[$gq��e.�����d�y�q�is+���V��_�$�L E���z��38^��m���?�L�<������Q��z�E�"x/Ymɔ��D��I����P2c��o��)�-�t��[�x�E�o�L؜W�%,o�����漾��}+o@� ��Ig���� I<9l�f{/�)�&/T;+�hc��A�(���tH�Oɱ`��k9F2����܏ ��?l"U�"Q^��������h�I�_� e�_���Qq8�O˚g�deS�Y6� �Gb#��NvDC*�$�Hz������?��`Ь*ADT��cQBj�:;�PpZ��1g�J�����K���E:ϒrJr���2�C�J�K�OuM�Ҭ77ש�v������)��2?q��m҃aQE�ގ�F+Y�Rm��'�Z�����l���w��$?��V�z�0���-0,�u�:�T<\O-��VHt��G��5�p�:�r��W/���@gV}�ut��Ÿ�����ֻ�{z�\*��O��4���ኍ'��{�	{�]P��&׆�uc����@��T
TIĦ����]wnm�r��i���ڥ�[�����.wO�]�A�
Q)���)�c
�,S�j�����g���iN���P9*�:Y{��X����(:�<��M�Z��l�PU�H�׏���7���v��> �Xx_��xy3�އE�eK��EwvF�6��꩎/�����[��8'����Ⱅ��&ԃR#o���֢�i�� M�S:����'��^��H��X��vH�ϧ�W����*�G5���"���*i9 ������O� ��k�qR'��r���\�xPR%��g����R�E�el���Q^�e �Vd^��_��\u ��m>�٦�8!b-�
�B�2U{�{��O��"�,09�t?f�ZI��������
�u'�ƿ�(ps�'N��Lv.Q�F��|悽j�瞕�(91lA�����+R�w�V҅�	"�oc}��^_eW��><|�1%�7Y�iE|�������Y�(�V�Y��O_�&v��f�΄�sh�V��4햏�P�.�y���D�	G�if�Ś��r�2�l�	�2-�A>���M�e�#=m$�* ��9����}dF�½��e�r�D�֫�ґ���	bq�d9t񥂈��������ˈ���᭓[<�5:j<�j����$�"10f��7d���u�D��}�@�gڅ��[݊��"�qU;��yÖ�|��{ 6f`/��Y)����̢���8���?�W���6�ɑ����V��y�+ə4�����X&��e�ڡ���i�-=5�i��%HH!�E��Cv&�do�nش�s#twu|��]����{�;KT'.��/Ԯ�Ǯm���H+��*��lg�%��t�e���CJ�����gYUsE�h6%ώ�k�R�`��`_������6
��#�1�0`�Ar�nw?�!ﾳ8.���o�J��7eťDv=�K���.h(Q/�^�J��)�hu�,� �^?������y�  ��p{���i
��/���E@�j:!����^¤�Q߯֏l7���t�C)�R���i�tk�b������敏�*�xh(��u��U]��1Q2)z�I����pB�m�E+��_��<�ۤ�����}�8�Q�]�=��*%~�؏'���5��R�r���.��;A�̎
0����[{���B�Y�A��� xs�����P�����(�h+T��~��h_�b�jZ�Kb��U.��Ewx���h�~�#�_��r�*/dL�����Y�2ܨ�od��v�����*���Qe��o�b$R-4q�P���W�^�'n���p�^[<_7��Ľ�TPW����u���)v�
�ț��;0��y˗x!�p�+,����JB~���!4�z�sW��z8�����s>�U��?��A7����m�����ㆀ���꠬TQ;WV����9͇Co���?��M��{+u�(\u���^�J�2�x犙˶N"�M��ү)^NI�.�s㲌��pwr�%��
R���w�8����`��;��]j�t�pT��_;�ؕ���������G(Y�wy�ď� ����ۚ�:�B8⛘#�h
��|�&í-����Q�U��zz��!2�O+CiE=ֿ$��%׈��m����`?�A����pDf�%��S/Z�e��*�E��3�Y��[K?^��c٥�7���t>3	�b϶���m0w{���U3��E����>�o6.W<R�N:�9:��R���+��.wD���,R���b�N'��I�	�f�	@Ɛ�������`�)�R�����֊�'յu�"�1Y�t).��3�+ڡwՎQC�m��{4Au��ۦ�%��M���p�m1˘�K�\���	fX�\���ɑBթ�4������6~�X�N���&LtmU���3��gHa���'Y�R���A��iF��� ���}�Z���t���i��}��-����l!�q����충��GV��e��I��Z[����"h�`Id���`���^(oC`0�</2D7���8M�'�����V�����I��h(�"X��s�l�����p�I8\�o<R��o���nj�aLl-�9�[=��<~H���<KS��+�w]�r��B��|ΖL�Oo�/���$?͕>�
�(�+m�'��\u�k##`
��>�$)���!��*�$���O%��m��a9(b��*�T����9{�l[W�e��^�c~�+�M<�B̺��pƠ����t�<�z��ZT�w[trp�gX�FD�4�G�4p�G�`��x�w�p%�f�]�����z�F��V�I9�|�3۰:��P�G�|V���[:��,�t]�W�;�fk����%��S����,X��s�A�ϒ�t^ٝ�$VX��[
Y���_#��.�p����C�N�G��5��i����n�bQ.�|X��8}�]�oo8�[[��!���S��Q*�'�=(�P��Z��)�j���f�3�s��O�R�*O�tZ����1G����. D�J�a0Y�*���v\�8;{<����w��kH$%�r��#�� �Z��ۇ��a@ �jl<�������D�%aۛLDs�����r���	%�P��Fۑ�:^������d�@�>����Ջ'�W���LG\��` �1�O�3��(DJ����x����f��f���=ɻ�p(T?����jg��zT���(y��{��8��� Gjp��3�H�!?�vv(��'Pm�iu��M`��4$����qƚl&��YF��B�kl�92Z�]�?vR��4�_C���aP �D���<��W�+��/�H��\�����D�??�"(�I�/��z'nx�$U!kC�ޒRE���qQ��D^��ۅ����?��N��C�=��S�m#1�����Z�Q�)� ��D��}N_�!;��������HE�;���=ڞ8UP#>�f	�9���HQ��D4�kkEu�n5)-�w��z֓F_S6��H�\��΅����i���K�e�3�+�� ��z�-K�H�r(���G��LδL]���Ͼ�2,�П��"7���z̫�<��d�hƻF1 ..B+�S�S��:f�����I�:1�D
P3�z���(b8��� ��&-D�\�&5���"-!��0C.����3y z��v�;]��QĶ�AWn�[�xs iVO�����!U�`
��N�:��Թ��Xm�\:��;|i��4B�|c���kʟ]#����qgq��fc6�����.�:ƱE��y6�v���l�G6&(�Ne�r?�������� `�^{��2J(�[�}����
��e����^y�V��7ϐ6R88���9�-�����y�4[�*�O�r�>�2��v�XO�&E�+i�u5��SXqZ�q�;b�<_S��&�lrW�E���O��HV�+�����!A/a>��7ʠx+��X\lG&�.�;�eY��$�I�X�Z�����M��C��;�l��(Z��)��~AC?T��Mw�}�|���G6ޠ2zU�i�� ����V�f�F �%�?�ؗ&y���(,J��8�;��"K9�I����lS=s0jMW
�mY�yT���;�E�3' 1{m�X�����JDY�3U&X�����kߕ*8�Ϥkeɠ%���
�� �5�r?*��І��,�ۜ@�������q]D�Z�Wnj�����LV���])��۝�N��[�XFEgTy[��b#����(W�����8%�U����h���4<�~Qy�����>0)2�y-��n������Qo)Л{���kp��+6�ὼ��R6�h6L[Mw"�S^'~H:���x=(w��߭=���h5R+�3eU���s�����x����_��Dw?�@&��/�T�g���B>�4��Sy�(��s�O��X��o��M��&d3�F���e��}��/Y��tCԀE���(�Z�)qR:����zwef`IS��x��+9���[�3��_�${�E�C�;&}A޴��Z?�A�1�D"j��,�
�jLr��F����;��_W��5#��Qu�'���C�;���m���kh�8?c��%����XhF��K[��Y�`S�:4UA��U�;~����
��X:�2'N�0�R!��s;�:��w����t�tGox&�G�n=.�bW�?XTC�u�f\Pw �YsO@��ں�'w��\���Jc@��}j�u�L��|_�!t��̼���=z[ߥ�e�CIW!�g���`� 7�zm�x��p2+��iN��>���CP��ݤ���7�B�0�q�_k�)p~�5}���ؗ���*�-�1	�;6��#߻��_F6��sYC�z��Yʔ�Mre�=|9�q��](+˂'���ZO�����w�9;d�k�c̻7��}��zH���7V4��N�'G*�����U*d`HD��zkP�V|��d��l��B������+m �6"`�J6��'���<�/M��=�)��i�@vf)�6�=H��� G���bKƇNv�ˁ�/%xA�g�
m]�f1c��I�&9#i�O����>O��e�^���H���,V
[�c�G.�����p�?Xmh��^���OF�4Ye��g�7e����G�↓T	��VI�}yغ�9�O[L���ۉ��t�F���G�3h;ɖ�Rq��J��Q�e�'g���/�Q|�*ɫ�"��ғ�4i��N|}�k�4�8-b�i�D�0�#��M��1��O��--��M���h���sV��+&�;ite ��"(�>�'Ǿ$Oi��,d�Zp{��d��ݠ�Uܹ�[o�_��H��Ld�G�E�]'�wvł�
Hq�ş���,߳w�cb��Ⰸ]�u�^g�ӆK�9����Z��4?6!i��~�$���$M�����%>��"4+z������5�E n���|,� QߺI
����h��4 (YW7���RA�L����1`�Q���Ŝ��lI��(�4���9��*p][�ҽ����`��D	F�9�����l�Ea�x=/
7�Z8��=[w�s�F�����8���z�|3*O Cp#H��7w�̙��7N
54�8tb(�'$���	>�c��vֻ�p����Iޟ�"1"�q4�7�x�(㉮A��ڻmE�E5?g�n�A&9�e{<i�.�\Xc���� ���Oq���{���pg�c��E~#'��h��˕�k���a�ﹹ�լ�Ӂ��ZҺ%���tO#��<��`�	���s|����I$i/-TF����C�X��A&��0�B�_�>��m���_�I�.O0�a�	��������Ep:_�;�Ţ���?�.�Y�l
l,g�5��8
٠Ҫ�C�"!�B�I2�Gn���������.�%q6Z��6�	�����r��a��Gi���Y�D�z�~VA<���W� ]�/�9���Qܹ�s[�"�#@��IS�r>��Ǌ_�q�Wo�<�WG�W�xj�x�m�<|>��Fb���18\���l�B@tI�CՃ��{���el!��G����Mײ�R
v�ս1���3?%�ϲ;�`�ٜ%@��D��1�V�!x;���R�q�����;J�����t94 �<�$8;�t�_�㚫�~��Z���~�{ûi��� �/Ԉ��"e�6�X.�7#�Ç�8�^��@�jjA@I2�L��0�Տ�S�%�B8��d�(�c�i��ĕȕjf����F'zUP��)f���x�I�Vd5z�~VЌ��5�O�\�YxV������1Ź�����5�0�2ЎI�q�)?�Ǯ�k�\C@�F���f'���S<�h����L��R�����EU0�5��B)\bl�Jn�o����|�� �cgi�Mn��T����^z�U��^�;�x2��v-�GP	��
M����_q�>deE\�ƒ0K���/�\(pp���|�_>0��LI��ꬍe���"��F�&
�>���t�Ǫ�1V?�hR�P?9�:�VԚv���h�u�������F!��1S�8�|{%���2t�cC����s�c��?��LP)˿�"�M��Jf������ح ��N�Z2�L�F�e���?����s�?Ҹ�#]y���(}�L�5�TЀ+S�Di���^֐�k�p\��.�EU�^�6�4��=r��	���rUBJ�e+�93�P8�#}��>]��D�� �Oιi��5k�n*�$h�J���B�H���Vȡ�}�J�;�]���s/���*�o������'_.Hu���r�� Or��Y���v�S��i����9��(��?��!����&6�E����K���np~=�'(��cu+���$,JK�z�P�sl#/.�w�rXx��IJ��ΟRisQ��{�GT4)�e^`�J�N�ʒgQ������[ Wj�,�3f{'��@Ƙ���B�%�`3�u	x�M,�놘]��&:��Jڏp�l}o�,>�����L�=����R
'[�H_9[YVo	��{�\��$~�`3}�y����ro�X���z�'�Bj�1�[T���������2R#���@	xcQ��*74�.�����U/#���� �vt^q���Op��7�r��b]YMX���}OD�G�r���Ӧ��j%��":������!��'��;�CJ*�f ;��DH}A=�uXM~Q�A!����9�3`4��en���
Z��]���rn�j�'�I�t���d�#��L�>;�;bMȥ.'!�+�_�/���O5M�^iX�U�27�	-�����5"%���-�Hu���27�?� ���S5Y��V�CB�v�L�-4��/=�`F^������-��qC��hDR�鐷ة8������ڊ|���e�A�9E*G[s,��P6��� *�T��f�N~�'�ZE���0�4!�E�.r��t����}��T�ب��vV���!p��b�7�8��n���Z��N|Jg/���9Q?ؙ���x�D��d��h��)�]���_b��=�W$}x�a�3{�4��Ր4v��A�oǇ%j*��Hȷ�t�ҙ5w&�2w{�7[����܆�	�aO:VrU�.�l��)<2���`v�e��e[�	a�LR�b���N��"2f5�y�f��ԕ�KMIu�w�r���3�U��T���ݔl��k+7�禃��p��{����&�'Ӵ�����P �|~vEr�0'y0�Qu@�7���g_���T�b���]�3���9jOHͶ��X?N]f���"C���`�Z�_*�Ȅ��P9�n��˳$��i;�h�~��S6�xir82����*a��0�n�a��Xć���F�2Y����y�g:���ċu��w��	hVD��@t�aat�>�o�]�y+�UbV?�$-�&�0`�Q^�e��g;q���0���4�_���4C�6Ñg�JB�p�t��q~���]���r5�kKv��i\�/­�%\�] ���:2:{��M~|��_>��X.P��T�K~3�s�.Y����9���	��D�|@aL���J��׹�s�Xţ��"�Yu;`��F�țK�?�� L0?�:�0����
��q�1���,���b�s�6!n�l�N��42�b�9�|��{��i��ு�peF������k�|�fA�(s��&VF���ܗ���|֩
[0��$A.��ti'DV	��JG-�
?�)�|�&��m�b2Խ�$�H��t{�TM�a���@�����=[�mHVT�j]�d��㖜�D5�=��+*���kY���t.)�0�Ya�U�"���D#�$���Hbc����{��X}0|�����}�W���~�����B!R�}������B�FauR"D�s�n�{��&�^�B�|���X�j���0��P��X���J��ҩ��M һC�]�T|�8����nȢf�T��i9� ��vIG	�.5r0uF��f�� J�Qk��0P��Q�̠}8������[e�J��S��F�V�Ŝ��G�O��pLԈ0/")x�,�#� t�I�W����+�͙�s,_R�k�ߩa[=�8��s�}bbX'ϡ[WI�A:�	|�+�*��UL,�ĥ�x�E)K3��iJ���v`����.�@�.A^Ԗ�?�Z�6��=aԵk�Ǒcq�M ��5~���AF�S���f��J:��*(������^����� �˕>9w/��^c���X�����N�-,Dk�Կ���L'
&����r�O(���o��#_ ���1ֲu�O�p�	�\��7(��"���g-���)���\� �qfj�����T�m��G#5m&�(����cjc���$���8�rdc���D{L���p��Wo��`
�d$/���1X(b�)c�n�)�!���d���??8{��������t1�yj{��k]	y(��M��`���n�z��Sĝ+H�g�S�Q��O�т͒�3�&�Nb�A��&6�`��g��k�Ynm7sc.�q�Ĳ�~��������ilW���B2�����<$r�sv��؞��T���y�o�
7�ߥ��#B�K�nͱ*7�[�0�Қz�;� ���b�(0�!��])�ϐ� �˸oy�JI����w=$}X�(J2�T��"���ywXX�G��jH.C����GBHx�Ex�D3�}��T�TG�Q�I���5ĺc�H�,�Kle5c���2 
<W�yJ,��ߍD�C�?Q�� <�!�)|��} �w� �3���!I�8\��ӱ{Y�T��3�OŜng�xI����èIb�m9��*zO���5a��e�Z�z�UO/o��H���'�$/�'��<L���ev�_��ī��^h�ܙ=� Nv&�K�5�*�������qfz'����o.���4{�\��ooK+�Q'qt�^�=Aϯ>�Ѭ��Z���I�c�����S̨�Ax���X����Ro{W���P&��Jhd#Ð^� �Z߼(�p�߸���0y�5�\ɝw�� ,��l�טۏ��x���&�j��UQ�N�%i�����x�������$��eP�[���$�V��~Xh�l��U9���5�,��0��\B�v�X"��JP�j=���ɕ�_�'{�b3����fF:>�
H��Y�G�Wd���PAk�(w�F�Fc}��W���Y�}�^w�W=���w�G��mg?"����jT�^?,����y�H��'���S���D��8�ʞN�]��	s� ]�����@#�����W~�lbB��{]����ܸ��0�,�{�פڐA�QT�� I�q��e��l�",���W��o�׵֭���g�Ƌ�����Ʉ�#+��µb[��7}�ϳ�G،����%���Ol�*�z��絍��$�R��m˒4v�`���G���sM�_=��mH�੒'n9��䖋oY�^�Z��^/Y:jl�m��)}��:�ՆAaW�iHc��5tE�#5�sz:�"6�\�:߅�9�"���w������z��I ���03�9��T�,w>�C�Y���S����"}`/�.l:��{�V������-	�mp������[~˼��"E��dK�:�/#%�
>���t��Ծ��~`��lAѫB����B�'��[x��H�Xr�炌q����#�������~F�1���;,���@u���Z���h��O0
n�����iᲔ����"�Q��d��Jn�vӊ��Uj�o�F�N�0�0s>��[�
�!1���X {������V!f���Q�얎�Z��`�^�aK�x�7�I�Uɍ�*=h�'i�U8�5�!�Dۯ�O�{
��x������ƴ�p>c�%�Hn�h�GX�n����&�����iA'�\�}���&Z�#�>��1�1ф�~��A��y|A�aEA�	aqr����oμ��Й��XV�ۣ�_�mf;�x$�iP��L����x>��&�`\��ʸ�bu7��Y�B+�`$pJ�p��U^�pX �ium��V��tOU�/8Rz�}ɗ����N��Ќ�⭥�q�b1�|u��݀��������')��X�\���q��&��3�f#%�eZvs%�%f���%�ݼf�+�m��2�^A�2��
|��ߙ~�KZq��_�V�.��o��Ѱߵ�/$�sH��~"�v�g&����1� OD�b2%zu�E�V�-����V�����\Z#&�Z��D D���"����Q�����BH��?�=�D��uJ�� ��#OÈ�v����U�>�Rb�k �h�wM�:��^y�o
�(]�?qhx����S�3��ƙ��<�D�g��gh�]Ԑ�`�f��6���{Y�s����?��Kk�k��ɥ�7�sׯ4�.g8B��c��Hbz�/`�GJ`j�2��FYrQ[��n�g(��X-�(,yE޹*WG+J�&�S"J���c�@3�.>(�@Y*���tb�N��F�񖄹R�����4Km�<�^�n񨵨P��%��3Ҕ]�����5ԍ�+��:�%�\9nŢPo�yf��,���C�=��1;3D�j�N���0����9i�s����p}���hU���\�i���	x�
���o�x�uӁԀ����iO����?N��e�L�ҝ�kb�CU�q�ۆj��-�ͥ=��݂�ȩ�^���<c��[��-!Q�"���������P��L�'�܆���܏ �^,��zX84��%�
��[��x�Mk!�♹���V��.nݔU<z@���l��!uo�Mo��2��@�������\� z`��R]G �����yz�������o!� �A�����Nc�[�J�:��_W(�Z��G<1�}n��[�� MG	��l�@�Q��;?6��	h2aE��2����MebĻ��l��KD7e��`.U�j�i����e[x�E�1�=����־�e߲�7s�E�c%,'���N�������(	�1/-�`%�F��+�)$x.�Ƴ�:�?��ɸi2��U��1p:��(�hA�F[
�F���9?0��ʿ߾*�e5�9�S/�>�7IIA�(��R9?�-��4$��Q'4	r���;�ˠy �Z����Cm�劰=����1��i�:^9�h�&�=�4�����0��B╹��w��*��ŵ�܇�^�τU��D>���Ƴ��w@1���D�E
�P^M��~SB0��5��ntP`�H�oZ�~�&���)ho����%����f|U�
7�W�6v�˾:-�:T��g�����4 H��	����߲���k�� 	D� N�P�]TDܲw�nD�\�UĹ�� ���)."�7R�N6�-D�sg�5k'8k�5n��b�S��)j��n���p��}UimK組>���)��%m���Л@[±��r��?��(��NX��l	Q�lZ�̩D�&�u��,}��r��AQ�sK��/�9̾�T��!Ӳǋ��3�9��̖�Vt^��sBn�:h���Ъ�A���	�2yMr��󰒊a���؄���/��S�#�Y�Ŗ�\@���.O,�5f����1��%���CU��c���N+w	ܻre}���r��ݽ��p��2+�A)w�s�As��gf�0`]R}�*�(jX���S�Y���	�|}�Cm�j%D	^��f(�j�b��8}�1Ŭ�^����	U�C���2qW�?gd�����qw�U��ike�|��.�`!p޽2|����3��@��k&$�ǿvl��+��Ne�������d��n�)�L����6�D�DH�5U����X@�<Y� &]�f�FT���%�N�~�t��OV��"Fvg���ib���62�w[�������ι0�|�q��u�ƀ��UZ-9IP�,��\:>�(Q�7\�7+�)"�ԏ��h��\�r��v]'�(r1}A�ʖ��J�MG Z	vT=�Y6�ٴ��,����)o7�n��q��CFJ���"�{�����+��z�2A�X���������I�n;g�o�^L
eDzq.�ų�f�
����&����o�;��0@d���l5X@������ ���P��t��5�������{5r=�,{UKmxՑx�	��y�*��`�����1����p�%�3	��A�0�tVY�E"�*%Z�4����D�1D�"�W�D*1�)�y�F��� ˀ��1T��n'�Gƽ;���^ew-7���w,�d�NjBi�_}PrU	ST�}���b���K� ��]�l�:�A�S���,� �[:�#����z֝��>4)yֲ�7}��;S��1�e<&|�Р�<�ZD�?��6�G|��/^��}��;p{��]�)TA�o��k����j��X`��	9�n�.�l��uD?��"��j��z<\���?��.Dy?����qSB�JIw�����*H��G����*��?Bg�CC`=LXmb�(`�Źp�.0��F��\�M��)U�pti�O�������k��~�GÔW�@f�<���m���c(c]�$'ՌEuג1�/K�0 R�v�����f�W�N�:����y�d�Qf�@Y����5��{�'4�dˍn�@G�?>?><Xl ,Q��`O����-�6��Q�k�eޡ��sM0
�\�����D5-��'�ɮp��Ä3����Zh��%������*���1e����3�ĆL5��6făy���F�!Cgx�P#�h��T1 ��Gsp�d�0���/�gK����ш=�hC�2�Uˣ�#�],>��?���@t:E���ˇY7���d�@�Ln.3���L�.䵈�&J��*�~���+f@pZ[ Т��n��Ɗ���ȗ{�'D�q�����E?��<�����p�'�+���?"�0T���C����O��c�M#H�l��؅�_�P��'�<����RJE���n�f+��r���
��� d3�JI3��U9h.���u�E��ABZ�Idֹӳ���`��p-(�z�S?��u�t���KQ1�"�G��ٚ�~j�qVZ��l�4�R�>�p�����E[�*�}M�y������%������؇�G��D�= �`�	�]Z�5w<�?�rHB��s�6�jz[l25^�Y�c�_H�'�#�S�v$ nN�����g�s�֫~:k͓bE�޿���~�.9�ǚ��!����hCv4����`��o�7�&'d�'�"��&�5$���ȥ7�T:�]g�]�k�ǨC
��Q*a�F��)�u�>ɧևh01�/a���`��z/�<pJ_,5窋(�â�ݛC��+����M(a�q�D%
���B��'�H��S����`_.1�@I&���妝�$}�$�\;��u��&�N�l�a6&���*[�+��2�G��3J���d�J�f�G�\[�c��#�����,:ySC��)�'p�t?����L�]�&�� ��E~���,@�n�z�i�L׉���FA��x�� ۰uE�p�{�i�1�Se�07po`a�nL9��e]�Q�),��^̤:D(:D̄��aڬ����U����o�|j����^��+J�nIa���h�����HbΚ@��z�᷵���8Ӈ��(��X�A�����?�݌jK���T��՞�2�U�4��z�Z��s#F�lZ!Ѧx���[AT��pX�J���*'�!̙���S��7��X>�5y���2O��6�=�ƞA��5*SV(�j��=�w��o���W���~M2����ã&a���A���h�$�17��q.���`�X5�A6D,_p�0�@)�V�,3OrAm	B�O3�G���8&��
�Ы��a"u�ӎW~�&4b��ac�Q��d�X��#pa���^���y�L����E�����4�0�!��?E9�3BR�[�y����ؒX���}h�q���Je�eKN������o��/+��c�8\"k^�h1Z�X>#�k���^ߔ�z�s�l��O۫��� 	�2��>�xY6�{�:E���/�^�����9���:����}�bD��&���b��c�~������h�4qQr������+�IX��@���%f~��lτ�&�J��L#?�Y�u�Y+q�+HB�5x�0�g�_(x������l�.f�c	Hܮ�<174a���4.�55�����t�����ot�\�g�]���XJ�+�E<��lbV���X��|��(���M�3*��uO#*�>�C�?��qX�q�-�LXR+���To�I��|M���A�O�q�e��4��%�0.����P]\��Ji߬︎�;��rw���ю�$� |m�U�z)4<���<�� ?�$(3rP�߆D4�p5R�����P�~|�)&�Ω��3ĀR�����J��;Gɇl8x6��:�{�����K�=�-�D��}����]#���DZm�y�M�[d��o�Wdh���d�
���=ۅӺ�/s(�)�[:�?���؃8�36w���CG��=�y�m���	�˿+-,���3g���iL_j�Û�qU&oKU�7~-�c��!O��`=O��I̧q����tѼ��[pr�2�W�j��&���osF5�:*� �B��OOO��B�S�V�'f�Ul�P@����{];��+~� +9�Z�gq�e�:�bp992ZB��#���t�wVA%����g��?0{H�1��B@���7��hU��A�6l�l�U�'�<7wy`�J����ݼ���=��H��w�z�r��.��"����딇)� ĝ<!p��3x�HlF��GǏ'7MG�މ)�b�u�A�� z%���՛��tPe}#�n,�pY�u�͹��d�V�����Ws5B0S{[(Tg䙿�ˮ�Hc,����R��Qe��W��Ӂ��ʕe�y|Z�g.�8�`�����DDhE�Ը��Sm�D�_m�Nz�X1�j��,�U��1fԎg�n*:��ش�:M�s-֛^b@E\@	~>y�@�P�|�E���4z�� b��Iы�A!�������KZ�Tki��P�� ��u\ꉤ-H:�)�>ɝy�^�Mv�|��`���֚$�U�Z`��#`桝.=�C��_�.Ob1
5pI�'T�jk�z�������e.�pU_=�P��Dh+�2�V��ǜ37;���Zx=�T��d�(�6��<\-`#c�^[��8N�R_��s:�_���0�'u�þ`��j��?����S��T�0w.VE�}��b�-���G�{�@q���D�y%���ʽ���MU9H��Y�Z}�rQ?����*���+��W5WW[4[@
�*�(r�q�n��2���i�*аے>:�$A	�#o�t�|c�Mz#�6�h�5&�1덩���R`C�U_o�k	<nշ�"�� ���㮾''F��N���u�����ԗ�؇��<(���7��o�D\���fN�k;86�[���A-uU����n�| 8b���P�;.��[�!��գ�w<�%�#�}��a���ᾙÜ4���v��c�ģ��gg��M!N��@O*fH�F�G
t�d�m_&��+km'�n�/S�d�g�!+?Bـ�.���I��깯��KNh���,�$/f�ڒC������ٯ��`S>I��3Rh��x#0�+�"/�����6@��ft�	,�W@*�dކ�gM�"��������k��]�O���r�/��P5�����:�mG8�������ă���4�q�����|�E���

����=)��zS�g
�l?N���@���"I֍n���EV����7̽Y�P�u����q;���/uM��o���P��I^�Y����<gڂ\?�$�Nˈ�޻��2�7���lah�d%��XYCֽ���.�$��f[�P�>#�O��* ��t�au *���t�.��{�~���	"^�5�y#�Y��@�z�Y��K�U���`��
l��[��`�o����i����D����pb6�E�b�*K���kۺt�������2��P���k�$gḑ$T��������Y*4��$��	��vֽz��F��15Z�"���tz�:a��8ȷ�Թ;���Bγ����t&&,1V�p��G�EJ5t�e�Єk]�����hOV~����8���� W��Y���/�l�>�q~�NJ�!����3)��܋��i�sz�:8��7�䉠0�����C�P��5�3��,vQ:�� ������ �)�����׃|��b1�_�?a�Q���m�-���[ �����O,%� �պ�C�����<�[�e�ۆV��GA��bms|ҧ�>����í�P�2�(SY����{�r����o�A>m�.~=V�C��<�H�6�3�{�>f��Q�X� �2��-�G�>�\�Snʈ�o��+�:�Z&x��TĊkn^q��P{0%�OB7��0��`;�Id������[NR�r9�R�Qy7A+հ��)�s��>��"\:<��3�a޶Z�0/�/�&�cO���Z����$�ol��.���i�^{��D�F�-b��C��Y1}eOvƐ��n����R�����[:��}u -�_������ O&Q�!��EXRz���_u�=�ĀJ�lR͔��H��ju�iMz�	�~s<�ڐ0��-8��
�w�2r��D"�`�'!O�F�(Q��O�js,�n���zu�q�׈��4$��I?���q�8���&r�i_d��}�n!�0�0�!�a�W咺�s�Ih������+g<
��жRo�>�P~��cNe��D>���'̡�s>� MD���vbI"�W�s+9��J�С�Ŵ���ĬI/�B4m�����_^��JØ�U!���"��+|?E72(�c���)E��$ow*��&qi1�gkB�:���R�q\V�V�0 ��x��qQ ����F���g��!Q��&�+�����S��
#�����y�G�"̲N"�yw(�\S�h̮k���r��7�oWG�8���v<\�3�]�bS֚A������x�D,2$<2#Ҹ�e+	��S���p��@�E;_���X�e��'��G��U3�J��f̪��'B:%9-0#&��89W�?V9���w �{o~�w⣣�T�/��A��Ң[�y�F�$mp�l�Ŵ�w�K*6pG��q���;��v�����[�&J���b3�eH{�S/̛&�m��51\�d�_�ڋ!:N�]�Z�T�߱<(��[�rsYY�g���:��	q�271��.,��H7 _��|�c�2��C�%ָ�F	ꉮP�V� ��(<�d�^�r$9��e)�)T�̩���R��Ad���=�������VH��XH�u<�ӽ�S*���
�1]�qn�2Ի�mB7���u���r]MQ������W"��W��М��tq�f����AAXie~$z�i��ԟY
BJ�P�l����x-�E.��`�X��QS��+C�B.u�o1-MW�Ǭs���@b2���8n[�)S6��7تR�O��[����m�9(���SG���u��1���'�p�ӝEŨ�d�?��(@y�����<57o�o���e	��8�h�_yK~����Pq�k@J3�д���d0�l^�ٻa����*e�8���]ՁV m���T$����m�%����)�v,^�+�P�Q�Ag���(�YeSlkT�brƱ���z@�8Z*���S���Oñrְ����PF�u&��c���0����|5�s`4����LIZ2;VՍ�=��J�Z�<}�P�~S�*Ƹç�^O�<�W|]L�!��ێ@O������;�d�K�-���e(�JMō�d���'�v�L������e[���@�l9����Y�{Le.��a7>��;5�	�/�-�(�u��UZp(4�X�{v����p�j�� ���Ӷ��
UD8�4�Ώ�+^jòڳ��ʪ=�\��,N�Y$^�Hd+�	s��&[����
������RM	|��֠��fl�*��OF��붂fJ�~Y`�{�8C��ƴ4��q�� Vk7�EO���.=�-�Ekj�l�����=��gr?��`�9���m'\ٽ��J���AMW�Wu�lz�+J�?�M	�|~��X�$z��u�� ��4^�����='�/�}���e�Ǐ�+<z3@�[�(Eb'	��K䱜�����,���`P(�n��n�x_�:x�p�`��1Ǻ�¤�ӳ��m����+"c���Q���-J�*Љ+~�ˠױ��� IVXx�#AK�B:vw�M�֯b]��$C��ҟgŋ,�#
���#5�X��k�x���GM_�2e��1��+�M��b���-���5�b>���=6)�B���� k����~� v�(�G���a��z]$Ye�^W�u��ۄq���D�!Ϳ�!|���_�e��w�;��"�� � ���3,WyW��� �:z�/�\�K��L-�'b}��:r�|-�4!dQdU�z���Vr��9�;nӧ��d����_��MD�?�q��	?W�˘�@�!���U�v�����
���X�ذ��[f"��p�*;�q2�cR�XZC�F^���E�Os�4���پ��q�Mm�]��M}��,=P�m���C�[F.h���f;KCa�S��/$u���!>C���BJ��L�kC�Y�,8���	0;xY����'��C[���Z�T��׆��Ϊ�"�Z_�`^M[P���˸�l��sY�8q���Iv�Q���q��-X0Cbz�����w�����V���;��xQ�<r�aw��C��G
e��*�rY!}�a�),%�j�Z����,%1�5ӛ�#�s�$��"�@2�@W}��J�g�f�s
�{���g5��@��Q�σ`�Yz��>mgj�� (*%NV��=jp�Nt�u	��هn)H������a�W�S ��M�|�c������9����U�5߾�W��
��F�7��p�e�e��F�5df+���t�݂�����9Ab���Щ�T']U�2S<
S�v��ɑNV�u�T	w(�A��i��]�&��b��q���A�	^ƒ��S���+�Q|e�yN h�P��פm�N����i16`Q�Sp=�1�k>pRN|Bh�g�A�4���ړ�ν]-R���nH��Ki��uln�sa������MeB�emv�6psū�B�����`������CƸL�>&I,_�".�>ԡ�u�wj��qm���>�k��
��	#��\7KH������Џg���_�3Q���A��{�	V� \xW^���%�_�G�5��](R~�:�@ܞ����U��(�Aݑ|sj�0��]ִm|p}BE�9RFs�Rϡ�j�c��=���O��I��W�d�<P���&G�N� U��|�&�粭�攛�h����!�]��pߚ�^,�.u(�#�4��0��%K#���`
��gd����Ok�1<?v�'T��vH�͔۰%#�����%h�9����@RwX�u\$�cSH;��D3ԑC�AwT��P�a^��
O����I����+(��|cɈ�.v�/����u�5Ĕ�E_�U4Ar^���*��^i�����b%��$�[�ي{��5�IE�b���ιL�i��W��wQ9T�/6CSyz��G��l�o�X���Ě�_(�G��lE}FJ`�ʣ�e�ئ5���
6�/l�8:��f�u�%3�E`6^Vz�gMط��}4��f�k���c�B��_���C4 B�� ��ŞT�~��Tw68ι3<ꌢ�B9�ߍ{8�U�K@��$��v�^�����]i&���-Y�ыX�0�* -�������b%�>A,���-:(�����s]�b �h����`٪�����6x�)z�����q�ҟ3��v�Gz�-���
2Y����>Q�n8L��Ԙ�<J71M�m4ߤ���'��@�N���&،I5�������rg����:6y=z�!v!� �#�:�Hs`ÈR}P�%�vտ���}�������F���Q��n��u)-\b��V䓤T�fƷ!��Q梥o�ŀ#w8���N�q3�nox��Czk���'{�4��B��� z�IL���<��-{A�ÆE�Z:��|v�+~o���g�Ħ���|��#���r2��~�  �C���=���H�#b��{ũ�����I���0���sr�Ӵ�K��o�Vxt�-�=�|h�F0��?�F�dL����l�C����NĦ�yF3µ����9�=��C�"��=�穘�����
�M�P�LеJ� �#�X'�qa�7	!*����8$
A����|�0��%����;8��d�8*`����s
[#'}N-q�?�(��{���Ҳ�c�� �J��"+D��bՔ�T8gҽX�Ѫ���FRc	��'���V��(󔦵o6� m����ks H��7xWa��%:�����ڄ��_��>5���^�!mO��ؙ՚�yw|��� �}������bt�r۶q{y�'Q�Idd�
�9�=�h��dƝ�ڤx������C�y�:K�)HY�6�w��?��y䘊�{'I�e9��;(/�L��Xd�wL�8Z��G7���z��:Ȭ=�ͯ-䇹���J�r& �Zd�+�a�x���׿n_u3�o��2a�G�:��G,�O��i�̮/ֶ(�ISLI��&J�f���8�ް��i#tbl;N5=����@[cŎ��zW�9�Dd�ΰ=��/�>�<f�S��ʪ�(��P3���!�|�!ke0<�ŲH
cxб�p4E��Ł����a/�t	���B��AϢ��Q#��F�� �v}	郞�(�1�L��o�����:����.we�/V�*�[�97Z��&+�%�j�X!�����!�;,�=�JwJ����0-�WB��:��1���	�!B�lM�4�ʩ�ee�sa?��*!6o������pg�~,�|#��T�26��h����E�9�囈��Z-Z���qu��[���J��7x�M�fy�<�>(n����MT&2��@?Xa�vJ�s��^N�Esք��f�LB�JM�U?�+З�8^�k �5,b?��3`��3��Q��6W�#���2��x���r�P"�5)y�,���P�E��-�����N��^�p��].��[Ľ�����`(:��NL�f�N�2��*��X�i�IF����a�V�+�=�Z�TR��݊O����1{P��5�ۄeҟk3��d�u�&������v�
�]"\��I��$�E?��x�kĆU�J�48����J~��UIa�ܥp�����7�;t$�78�D�*`v#�Y��o�Tr��y��RZ�Fa��L(�-c @ˢ��C=�i���N�`�L\���
��Tfm�x}f����
� �̏?%��������g�D8x�&[n%�)�q�!�2��x�SY��<�=D��&'[��6I=���Ф��|�S�H�y�<�����l z��������,흲��1�󺠦�*2U
D��Fcּĝ+�'�1|�uGW:�lr��et�o��*z��H�:QPW�WuAz�y��YASa�������f�E��]u$џ�����7,4>�ϧ��\�X�f�ޡ�J�<�������a�"�iEl�l�p��UMi'�2zC������u�L^Y{0�E��if�ԏ,kD�S)1ƌj�L���V��۲�u.Na����MH�IO0�VՃpCT1~�73�1�yhm����p��
���'jzjyv�À/�-u6�a�h`Ra�?u���K$\˯�I�v�2�»�^���v8�a���V���LK��VˊV���9�"���wM���e!��3��O���\�b�ח]`"�ɑ]r�0�w|�B�G��%�	�����P�xA��m��ئ2��t��A��7ۢ-Ӛ����!i����Cڀ$FS���9Zw�<Q��db��ټnꕛ^�z(M������;K(tY��Zz�=�˾�"s���W�<��R��Ȇ����0A1��ۑB2I,�P�����3b�������I�_z�6޸nZf�&�F����#dW�S�T4��}d���JQmw[ y�9�����h< ����O�_���Z=�R�P
�9��s������z��Q5=��iZ�Ѹi׽�`���o��#��FN�=�-�������_���H"?���`\�*Qٷ( �(.��P������݌��Vm!��`�h����lq�&0BnC��쨶mké���"�F^>�<J#����%0�Ǣ�YQ�])�X���������+
�%���6q��8&�Y���5��3ݽ[� �����m�.�D�\���X`dM�DZ���-��7�ėIuuO�#y@��.��X?Bx���o�c�^��5�Uƫ�G����Ӂ H�+�,Ĉv5j�_5��Tc�a{�/s_��Z5y{�;�<SOB��Fʪ�H���\�{.+��{��_SD���Z��5��u�.X d@�|��b!�⁭��"����;�p���v�1rGd�C8
A�H�e\1�����Z�:�&!hI�6�T �{G{~Y*�mQ��a���"��V�O)�<�k��2"��%�^U>�U�֊�x��	�X���"��G�����O |O�g\~����_��r����w�g�n4�Z�Xs�Ȫe߭���q�����C)���%���a̼.����!�!d	��9�A�@�g���Up�DV�N��� C�I�z��4d+��PzDUK�p�	�7ݘ��1>��a@MDoK����9�L�M���ʚ���@ʒ����hٜ4�9�i#��B�~oCJHT]v�լ5e�R)�Cͣ������D����]T X����:l��b����\I�F���5y�J��uɄ�U����X1/aKY���#���%��7�\�.�H������V�F^�����-`�aނ��RA���"�n_q�^,,��3RA�ȶ;�6�t�ZΫ7彂�,����d�
������s�.i:ќ]/��s���O�\p��ͨ�2���ޜ�Z��ܿ'�G�kT�8"c�z�t��Tp�� ;�&�! �?/�(z�Я�@<�Ͱn�k衫ٜ#�:�(������<�4%���Du�Bľ���I�Mðt�ض���#�d8-�vC�{��{�^�Ζ>p9A��~��	�NXHo���fM���=#'%O9Z<��,�AsEy�W�z�J��t=�c֋-�J6ma�E*%�����mrE��G�� IqDn;�� ���O������w��F�~$��)����
���z�f%��߁�)3�G���a]�k�hN!��-�]�wl���d�Ej�ˀ�W��Y��(g*�<W ��0j�"dQ�Z�;��"��ps�_�ƾ!�u(����� 4i	�o�9m"{��G/b� �	|p�gX����c���߿,�)F;!�I,4+߁�{��T��92���&Ր]�
���J�H���: �,ۅ+�_P��a-EL�0;����t�1<av������W�319�U.��_0�wԨ`Б�G�n�,�F��n&���+�7IB�ĝ�I���+��U�Oqw��'}���f��}/Q��ʚ����+u�u�j��	h�xţ���@.y���y�
�瓷���*0EƖ��[-8��;'']�{Ȏ}� �^���%��&!�R�)'���a /0P��>]��[��l	�~���������$�~�0ӈk�h�G��'iɆ�S@N^W1�z̢�.Z��oV�Q�VD��n[O�(� �Y�E��G1��j3�#3K,�妌�ཻ7=lض���4H�v�>�Ky�"�kL�e�wb;Z�~����9WJ��&����C�Ϟ���S���V�3��V��]h�7R�h,ōtZ�Mn*��ƍ5��N����.���C�\�@��s���$޻�ydy�t�����[���D��T0�@3s�+Jb&Pg��6��\j(���IMӀ������@x�u�Tҕ�ůS��`��jI[�+Ǻ����=����~᭙�充�Ϧ�S�
}a���{�:y"�vV�TB������a1��7G�O�%_=�K�C�b��MP�����?�%i�[� ���j@g5i|��%����I!:��s"�h2��΄1�-����'�%�%=7�������4�*�O�2c�x������i�64H���pT�fQ$�Z���4S����Wl�`�-�*b���\b^����MT�����t3]�R
X��].��l�$�gy���ol�����#^��6����kЀg�m��R�ݒ���v����^���{hܕ���~r�Ks�����9UJŏ,<�w��0�M��3��Ɯ��9����ũt��Ak��lS�%��o��G��;�?=��y7�d�_������h���5ʙ3��,;�������<���,wa�J�����J��YF�������=7���W㰳 y��D7
v�0IY*��]�r�B�QH�[��ExNf�Q�:Eѕ��&�Y������=Y�}����0��j*R(��A�J�"��wk�TJ�)@1� ����O՚�0��ݑR�U6�k
�S�ޔ��-����FE}8��7uE	7��V�;��^>^c�t1�2uuf�ZH�W�*��0�mLn&�G�L��O�"��m���&�� GXG�h*���v����	wyQn̶���/֫n��q��{��u
PaS*?��>΋���-R�@raVh��5��Z$w�ڑg�=����y��;[R=��@ĸ��Ef�Z�/�{���%�O@��Mla�lh���^��t��V|�@�����>���LE0E(;&wR��CR��DE��̆�2�;�
FT
�A��G��p7�_�v��Wu��cE�sqʬX�-��C��X	t���̰Y�,0H������~>�b��z��~="'P�p��g���¢�G.���>���
s���|��wP��g�ڻ&Ai�É��{�q�z_+74 �"��|��yD�	ܩ=��$2��I[G�T�DYp,=ɹ�$� T{T!�Ħ2�}�h����l �u����4TiM-`a��\Q�Y��\t���wk!��۟��MDg���O���� �߸�%39*�D?S����5�-W<f#�#��^qQ ��yNJ� �����"�m	$��6�;�m�����@s���,�Q�W�����`��+����T\�tMCTC����J��JYq�a�q�lsu���:j��9����J�
��Ȣ�ee�.u�Z�*�(ޕ�n������bJ,�#�GPl|1T���r�돭n��~��yL�@��B����+b��w�=���L�&�0�Xꮡ���ѵ��� GG��	�˽b'#k�'�J=ч��1ѳ�� ���<�.�����^�)!|�k����T��E�$��+��h36��������Kx_�`EV���q�,���C�X@�5Q?����=�|���VD�j�ؖ?��Uq�a2������a�UI�s��P&=��9.hg@��}u?�t��2��Z�/�ޒXQ84���D^�3����Jm:�I-���	){�<�5>��+����B��8��0h��z �-v�q_S�a�Hz?��"��̿!춦��9��s����=Ӗ*o�P0�:0y�!|IQK*�X�PtzL�����5�S���p%��v�Y��ܔ�O=�����Z��'t�����SH�Z�e��MIi��~o�MÎ�~R.kf�SZ~g��]Qt!5K���ML5�92��\JB&O�����x��^X|28�H�`i$kX�,�J�&�g,����X���i�-/]ŗ�������:u��4A�� d�_�9�R�����_��C���ֳվ�@�
ؙ��';Y�B����R�(���;*���CQ�2�\+�W�	au�Q]����z�T�~ʲ��E6ۮsq�>h<�|���E�ST���I�!l�0G�8�4k�Tê�
�)^�rd�؃XHsN,�Y+VY���^����E��Z�-$�t���	������	S�&ﰨ�/O�Dn����=�a�?oaF{S�O��hfwb}p��\��lDf��E �*͞6km�{"����f��PE7V�E6�A.��\7ˍ%jcfB���x����q3Č��/�jM�
	�|�W�"���)s�_��� kOэ�	@���͟��,r\�ң6�|��$c�op#�!mY���E`�j�0��6=" �޺�eо���\�%ӧ�i��a�����IxѶ6��-���Y�]���a6�$i�� 3�UX�x́�����f���m#�]���rԻ4א=�-4I��.�۷<�v�Puq]�ٽ�J�:~�{���
����,*W�V--ސ>I2�nX�X�(�8�ޘ2.8�d�ø-�]��G�k�<��������s'�R������W�2�'���\�q�e:�x};(�����@;^�����肩�Ul��b���y�G`Ӥ���R��8�X�k�j}_ά������fyg�@��ޡ�%{;������J�H��D���~d��1׿��Xb���G�J6�[�#x�Y��$Te�AK��L���W������qG��	Y�w����֜�U��C{�y]�-oG4��]x��5M�Q�t��{^�7�yf�18������ 8�cx�DaRS�p��zm�*9���%�B����2f����%�o�����{�l�J��(4:��Cs�v��o ]�����vf�%&�Y]���B-?=0+��7�+Ԕ#wzN����tnݶ4��.ܮ͜lo��*�:�r%&�~�)�%�}2�+Q��b�-ق�@j�l/GyU��*r��J�:#��^�Ys��X��|������C��*�e&dj��ͪ�li�\"V&��V�w�,T��U�y�	�(�r��8�sa��C�>�>��뺚|�"������T
_�q5���s昹i2��0֦�	��AP=��&��&ֱϫ��iM=�qʣ|��WW*��z�K��2��W E��,�S"b�E��Q<�� E�JL�j�ڒ���oi�XO��OSsX>�J+�wH�\_%n�C�H��(�ʑSr��h3@�f.��m⩡u�_I쥎�V��0�(�8IM�2���B�yM@̩��4�G��S�ӟ�����I�B4������Ȃu-����`�x�l?+R��ېf0�ܳ/Jc�Ka�&q<�"�2M m�6�]' �F.� 0��E��v��`�/zf�P��H)���Y;@8��FS��}
���2NO�BS@�]k�m^ވl������Q-������o����m6χ������J�&�nLI������{L��#l$��{KYGw��W��S֡�f���%@b@f�� �!t߮D/�d�&��ꋮ��@��8��@���'R�"7���F���}�:X`��pKӡJ��^AG_�G�y5g����ِ�ά���������?X9�^5#,�`+�h0�g�ʴ���I#�u��2��HY����MK�6����N�n�'�/���YG��Y.t5)u� ������+�{Ð�%[���m��ɖ�)E�:��K���6���or�w���V5�Ȑtd�s�q�#D���C=��=[����Z$��ty���;����>�*�&"q@"��f�0�#��}ٱ{^m��>��g��������z�̫57 �&�W1'6K��╊���~�@;���Y(�����s�k �]�+x!���烥�d�&ƩY�>�ݓd�)�T@l�V�� *��5�v��up[�}�#
�v�j4��f�լK������+ϰ[��	>�N2<������@@p�C�i`�w�C��i9�RK'���=e">{7{���ޖ��)%ɟ�ɲ��B�D���_�^�AU�n�}�V�Xe��#s'��%�DL�*i>���Ní�v	�s�1/�թ���Ҵ�p�{݃��Rư>�g���t��|��SA��Z�Y�&j-��U%`�o��5����N�ׄ�d�}s�;�uXo�?P�tdv�ڇ���Q���{����4CK�/�b�� Eb����~��~���&��v�?4b��Vp�'�0;�0L����#KCe����c)SiEV_Y�c�5�w��G����h�v
�Gv�;�І|#_�$���_�Bzocte)\U�B@�L��p�SL��)B�-��D�ܶqcF�a���/~�����h�^�T���l	Â3�J��&Nx��7S�ZD�dLR�2��zA,-B��ٹ�Tɗ��
ܙ�V���Tp�z�NKD������E���3`.s�K�0׎��2���oh��HL�R��+܈5�T�#]��#�9\X5���,��~���r�	2�G�t�ʶ��� !��ś��S��HH.8M�p�t��wΰF$���x"�
hJ�WU�G�Czz9��L���y3GkvQ5��8���JW���n>J�o�g;��NV��m�-�ff�K�zkr�z����T�P�n52f� O�Q�\y�6���_�V��=G'0��-���8</�9k�LX��e�W����<�QaH�Nd�����a20�`��tsv͞��P���v�$w����s��S{�T�p��HT�h.�L��åR�"/d�h�h����յ߸;�VU�m��Xz�]\�����N�?U����YYW�D]�]ȍTdH�l�=c�ݔ������;�p+eP⾈qv(<v񉭨�w+�>&g�k������տ�4T��!L�Xx�V�[\��[��9S�1���_��9�I@!����B��yl��͚���뮛>�kΖ7:~���<e;�K�c+Ӟ{[W���gb���GV�Gr>X1�~<�c�����l��yO��yϛF�t稔�O���ң��D�����f]���2��dܑ��������h���Ȇ@|�P]G�N�0ʦ�r:�8���ha�؞!�ӗ��t�D���g�x�d_��/AÜ��b��ehļ^�}/��ہv N�y3�X�;D�|@�h��K`���d�:����X����2"�M��=�1�� �E�t�7�c��>�i��m�H����_̔��U�z� ����B�)���Z��?�P�)���P	�n�����d-�hÎ���ت�uL�w.�����o��3y]s��U��劺�?|��!.i�ԸeP=w�ۿ)@S�#R�Y������7c¥$�l�T��)��(�)�#<<���
�yT�{"��t�u�&�V(�xY$�u}�����j�l�c!��S����n��At�����x@���+ʱrl��me���&ϢI<�a7.��FE�-+/A�pzE� k�m4H�����/ �Q'|s��3vj����W�W�:f�ˈ�<��-H𕸏���ȑ�BK��HɆ2И�	>V.�(Ut
Qr���D�ޠda���HO C��f%��*L0��8��#�f����`0�Vqb��m3%ibiKA�8���Ԫ�6��H��8\qG����<�	q>6Ws{ oh?�X�g:eo�c��py��X�{�^�Fg:�x���5�݇w� ��*c�rJ��w@,H�����7B�{����X����U�I�f(�4��7�	w�az��/eQb���
<�c��eS�i@&v ���|�/�'N\-��d��逅����v���C������y#�֎Gk���,���"�	��v�v���W�x�oљ�S�^���P�a7�o��D�&���
6&:k1���/+/'�q2(\W���+Z��T�r����n�a���Er�%I�<���5-�PEKV���1�Ih����+|�p����!����B_�����Q�1Y�$�~�"5v�z�s�5�Y��S�RYYQ�6�F�a�TRw��!����~�(�A��ؼl��.�ח���ARې=q�ɨ�=�>"�\������	^%H�*�ˌ�:�,�i'�D~��iNnO���E���R�2��&�ZE����ڬ�5�S��^u���'�U��x:�M���}4���U��=ع4������w�.Y$RzQ��.9(ͮ�o�T;�C�񇷂��D~~(J�~����̋U֢A-������A���g�E�Q~U�pC�E�AJx��z�O�����<C�g�$���V��mn� �����j��7mc��1�0����g�d�� �>�d.��f�-�b�����.����`�yR�oU��3���!(�9����׿���
)����)}u P�����G�g1�ܱsYe�Qv.�-�g�h��r7;��N+g�p[AP��ݻ�vpT$Лmp=XWqF��H����I�*��>�KIڰa����a�{�Z������(��e��c�dK8�?R���H)��W:����������C�z8��20�!tg�"���T5h��F_��A�k��W~�|�	*i�q$�7�m�L`�ܹ�y�ٿ��82&U�U�K�����vx�+9,��K��}��f^!��#l��[�<<��f?vk�TQZ&�>vp��Z[�XWF�Ho^�tJ~x�Fb�6O<-&�K��>�g�	d�K�J<� ��rq�p*�T�<��x� =��h���RV����6��ǂP�O�'��t*˂��|y�<`ۙU��+?����dϹW�}����ܥ�ciNhg�E���¦���S��4f~mat�8�N!o92��{1�.�bYo!:7�rO�������d��i��ʣC�X.�TV{����y�D����Y��wb`������X
<N���q��Sc�O��#Ɠ
έA��g��������Qcu�w7�!�M������o��C�!��ܼ:#�r����(`]2�,Ѻ]���V� ��]]��|F���W�(Z�)]]��}D�}��Wc�����
��9���ܘ�pbr�T���Y��d�v�XǕ��h�q@�����n��7`���Q�X�-cI`"�3� l䉹
���7�ꅳ�U���v���J�c��W��/y��4��O׎n=|L�|-% ova�ʄ |&�I����JT��Z�x���w��j�����Ua ��D��@����^A	�l�Qj�g�Y��kꖫw�G�	������*����=\����F�K*�j��/���[�u��I���YR�A�&B���a@7UAOr�*�m�� eŪ�!׶9�*D�3xA_@(_9뢺��~2�q���H"��w��؍��	��b�h�NC�l;ܒ�s��T���үpR:1�x�"A�K���c����LZz=D�<M�F�t�Pa�;GAf����b�h8��tOFNL/������lՊ���a��c��rg�l�imjsK��߮zA����ɴBo.ݚ�&�(�@05Ts�
��i �Ǧ�M,���!����%$7����#����w����b��~�1Lc쥃�i*���-a�ͧh_�c�I�]���?B<�Q���V��E `����?t���P7���pMO�[�������uU�Bmŀ�7�:��QƴNϗ *T�l� ���C�r����x���|Xk���W�K��3H���LY�v�O�d�g�m��&�Tv(;�f�?��5cS�J����r�_f����{�<�n����#���LD$�Q��E��Ї%C>�W)�����ϵ�l�,B˴i��o��^T�S�	/�ޣ�[^�D�ꪚn�w�u��~hT��K��D){L7�~��i��f�pARdQ�1�ѥ�3~�!�a��a��"J{!�gg)	QqmLf(�%��aM�;�v�v+feR�Gi1��܁Ü�L���ݨ�����|�_}�2kĘ�lukb.��X<���i$��������Jz0+|
~��\M�l5OM֟�����/l�&�b�V��{�!����=C�12�Gm+�Zڑ�Q�=�E:,�����p��=�\�{�^so��`�L���(9
D�w�J Oyp��Ù堹�E���dR��T`���\o�ܯ�$H��(��!e�	O���©�.�;� ��w�aV�Ɣkb"�Í/��f5�a�A9���C�;��~}�(f�<Z�EM�-C�{�4��5a��/�a�[@��z�����'�Y�1�-���v|7�M�C�t�P���/��l�1����Ha�ru��9k��?�4��u�j�c���q\�:��л�%J��I�m�!�����<ȭoB�=Yߴ�N�n�}=���%���-�g�y���3	]5��Td�Ϧ��kݗ�=~�PlA����S�g �u�^a�ۅd�&�榾@�����z��s�ɭ���q?1��X�`�~nVT��p�y�t��(�ŏ(V��3<�
ƍf�<��	���q^��(�ϑX	� ry�+�h��[~���Q�4�X� |�$��~�D�O����ޜm���_U��������{=�F��� O�p��U=�UEh���1:!o��݈�Ob�)�!�ME��;���Յ��zm�1癦�$r��y��T��ќ4���c+}|1�![�ʡ}�(k����)��Zb:�-��X쏂���E�_f4�4�VK_��I�N���M�X^o��=B�똊񞲲<���:`ad�b�2�qa�|�C��2΁f͆��U������)͝��p�#a���F�y�p�g������=p/���8�5gI@�l ͢T.����k�3B�}��t���G��_m}y��Puۅ�f,��j���lc� +���-U�T��-F?��_;�x�wA�C���O�x�����u#�Avd��Dx���ǚlw.����Q��iT��o�	oGv��[\�������g��m����Z����L�\/}_�.�����6��KS�(R�e���9��q��o��?����~Ry�]p�d0���ܮO"oF����@W��Qv� A�M�v$G�m��3������)�q�!o���Xߑ�ɈX.�7h(&���M�r�g;�$c�שm�sڢ*C^ԇ���2b9<�!���k������!���0>�t�(��b���i�� �_��(�Pղ��!�jù�C��5e{P&ȕ`�R?%-�r(<��'�b�l�\n,g������:�t�X)�;<�"�]㐾/p<���Rh0��j��Q6=�2���"d�a�-��f��y�/��}��ik��"����R>`�Z����i�d��v\ogVQ ��D����@%� S+��<���Ѩbv�2��n�Im��[!G=��$-�+l����!	��ԟ����Ŕ���?�׏9��E��$��E�K��	|'�v+�/���h��v�E�i����k_/����X������v"�����6���#C=�O����C�."E���'��= *�5�7�sf�6*O ��i+�)�J���Ȧ~O�E����UaŻ���O��>�-ZN�Pz��c���ٺ���w��i��\�!�܄�_�η���&��g&P�� �;6�a�9��'��|�}֞I��q*��3�x*���ܱD]��_�����xul١�ٯ�V����.�n(�q*�kV:�i�
,�W^�("\�� [����@��N>��|��Ʉo?L�AS�� 4s�\�3
q�4�S%�a���T�l��kB���ur�Œ�x!ޗ�͗�'�L7��7B�l=cx���� ��^�/���^�9/��!	jf����Yr3�m�
$�A��بM9 )�B�vq�-��p�0�4��A�@K��}A᩽r�_�屪�(���ezj|����q�	b6u�A�X �*�I�:��R�Պ!��)j�8�mJF�Yԓ�0׿z�e�X�JD/�'B�p�]�C������ �u�/��o��%��nl!HA'���z�p�.�\;W��F6��Nr=V2��a��>����h�[E�[|e��3K/�C Z�.�\����E��b
��}+o�K�u��ϩl�@g�����>ƅ�BɄ57���.�@B#������ �*�?Jv��6��U�wPhPkzzJo�|j���}�o�pv����?�]*�����k��ҽ#�xS�G�PQ }g��U�Gf^�8R �/�=������sn
71�����@��2?c�ځ_�N�����29�����JuLc�7x"�$qz����,��b�=��sG~��Ê��k��S��u9^Q� �Y�0$����pK�'������F^�_E��X&�R5��
�sz�9AB�,!���[	�(�D���N�Ɉ����$��$ώ�S#��/l���W��n~]�3�V$�L��evR�G`���R� &��zɫ�䐠m�n|^����J3�X�4C��W~C��X��N=���ÿ~�m���P�a��ϴ:Y"f��LO�(�v8�&��E%h����6Y^朢:�4��+7�B�~^ݳ��$m�{M��\���P���i`��辧�*�j��k�& c-@R�/�P�ƏP��/��r��ʴ^��9(�[�N������Ȋ4
��j��m ��t�����L���q�(&���`�ق�Z�(^�b�d࣪r�̍������cPi�;W,[�}
AAp{���wwt#Do�:OdfU�ܲ�oœ1L�������j��a[�Re��b#Y'ǹ���l	���xK�+K���E� ���Ο~���'��4rlz�+�*9�.�N�Emç�i������q��~��P9(�&f��T�
�\b��9�x�c�Q�tT�D��n%��2,�����@�e�P&��F��C�M��l��>>����wYu( |w��F��ˮ��:��0�|@�)ZFB��<������4�I����:EVwn~��=�1�����S�3�O!&P�s�_��R!T"���#�*��)T���p�+��O�J)\�0��v�ݓ_��B��u�o"�Cͅ�YC���O�:�iGq����?�V��oH*Ӄ/ه5�m��YO����D��@��%6E��=��O{�9x[���>�\���"(X�m���4KJ��(�ƿO���(��j(Ea<g�gx��:�(��~�|v��2	{������~l<?��N��l�OT"+�&J�a.���~?}j�]�Jݩ8~5����ޔZ�!���$�a�<Z)u}e�1�LT͜LԢ<
���mٙ
3��_�?�_g�;5�^�?���r��=��ÔcD/3=��l2���� 1�؏��6�*���T{NѪ$o�&<���]��C����2��
-Px����4�83�
P�
��x�7�L�Ҕh�l���"����M�tՀP��=n&�K��)"ǂJv�@�90b[
��z��5��Ő������d�!�I��(�;�]���zO��{���-ք?����� S��2؍� 鬴H�W���~N�'X�ݬ��D��<�4��t��6�Ga��ݘ��Co�݇� �?�Ƹ��MҳΜ���h��l�<��d��y�a<����	���KX���-7�2�ݴćY���ƈ�;Y��`�S"t����Ҿ���(��R3D;A2�a	�M�#i��%��%2?���6WUH�P!�8
�ꢷ�0y�T[��H�r���@o����x�6�lUI���>�L��0C,�B2��=����������,�?�����z�E��-���l�̥NjP�b�-��Ni*�Ay]�xgr�������nᥚ�d�����h���[�f�&���U;V貚鴴��[);))M�I?!,M��I������m�08�j-���.��s`�����a9�ϯv������Ն,W��=��(����u��jr��|����:*a
(@e�)'(]h�f�BnK�O��<z��䈆�v�څ���V�l�ღ��.n�Q6�r�T�1AuE���(sioE�i"9;RË5��]�Da���j����B��GCy�#a����� k���r�I�1r�*�:7@x&�@^t��孫╍C�O�7��=������
(.��Qv�A��a�v8}�͡�nhl��5�!c��Tu;��d��ԁkU�B�QAz|�TƐ1��U;D���xzt��^���.^Bf�;,��D�v`�ŕ�dHB�X��sS�v��pAAA��K�peF�j�N�����������F#d��~з�6�V��f�G2�,|KH�&�F8�Q��o����ՐAT�taXc�=9Kʸ�2��j,fy_[��HoAV�}��Q�>����)3	�i��=���ʹW��l��Q���BC\Z�����^tEG��wU�F[�
���8��V�=�\�V�5���Q���+�&���cid�E��@���>#��n1�_|������F3�_J(J���v�a�P��i�s�
*�ֽ�,F�%k�4vm�̈́��F2K��.�Ѹ�W�ř��P�P����D�P�ɛR��_q	�[ɝ<��6!�6�� 3���R+�1ux�eԤ���@lyD�|s����n�bzI�쯦�x�nz0�j{��!Ny�g�<Sg���8�/7����b�T��G/~�2Kۅ��Qp�Cl��SP�v�*��@t�sh#*/I#t8�s��(�V����C%_�^4����Gs$�l6B`"c�m)U f�*	e��.O�&f��.6*�{\���˲�A��q��w*�f���<QYiJh�8�[)��V����0�p;���k�� }�-:yu���������IT-W���NT/s�]�b��B��{)	'ffkfA'�z��4�f�wiQP9��SS�Ȫ�i.l�r�üc��D�(���P�f���'�[ld���m���#��ul]n��6U��b=B�U��1�U�7q�<�t��G�N�
}䔎�ł�ϑ��Ѝw�3��լrX�J�Qeo-5e��Q�t�M��J�D *��@�I?������MX�x�����K��G�>b���ZF�nG�~�T�g�Qm�`S|n}��E3�Oy�Q�w(��S��.���Ѽ�_�Il��v7ࡣ��q��f�B�6�rō��� �P����&��u�g�Ϝ���BH#�d]��s]+9o^�p��#춹�{���W��)K�b!j-�R�n�j���0Y/-��E00l�1��T������3_o�A�V��A���
���v�:�n37ݫ��w�[Y�����ƀ������@ȅ�2;���H$۟�?�^Z���9�; 5��2
�\ZV_����#P�ԟ�H�-PT�-�܂L�~w��H"7��Q �Q�d�#��)V�ܳ��Ҙ�l��)�Nj������`��N���G���T��Ɋ�egt���s#Y[p� b�Q�T`a[�������&�Sn1�;�&sc��
2��U�Y-��Ч�Z�3�H�~h#�ڝ����=sU�����Ԭ^)��_J>��9=޼±k,21�$pV�GҴ���}���Aۇ�T�� ���<U���ՠn>�ZÙY�ڥRt���V�#AH웲��my��+���g��w؄�4�d���4ݳ�^�zf�}��d�բ����h"�Iל0!i����+V�݈��X+�o]B=���p�B�%��>���������<��h��B7ۻACLnxڗ��1��n�#�1C�Ҧ���(еȲ��<d@����Ԯ,��s�/�ۧ�Y��6��ʤ��3agb�^�Bzվ�����p����$���2�'�h�����[�<2�Q_�R��szM2���Du�*r�٦��|W]�����و-+Y�%:.bS����'"��x@����c���Ϲ�@�X�@f���옖}-굠�����m���sY������?/��[���Ӝ�����؋|�>!����9	{�YQ��JN��yM���R�m�~�fL�$?Y�<ڝ��.��0�z�\3)W���#�T�4���"�7=Ə2}	�[z�8i���FO �u�[�a Uk�/�s]c���\(9��p@�=���bS�(�v)�k]�K��KiL��<*d@z��rfz��6����I0
;��d��P[�e�O����F�emH��P�F ͯ�=;ݑ
Տ�4`QW��;װ[rxX18�czAD�=��K�NvĎ�r
z��0�؝Ӆ� ��n��|{OW`^��We��,"���?�.�c��3����*�@��k��Y��Y��:�(r�������iN�$���r�e�f��!%*��N��M��~v�]a*]���'e�zq��ҝ�!�Ln)b��� P��[���V�_�:�N��m'�9��I���F��E���Q��O�q�̶���D���L�����)�����@;+�$�o-{m$r�a�Z_K����4��wX��&��G~X�.��ύN�0��{��w$�-�
��`��kZp3���"i�ѱ@�R�S|�Z(kCc�筩�&�c8`i���S�F�0��������ѩ�R��m5��{�)��y��؟я����6Y���k��T�@�m�o'�����tkdA�t5�g��`76[ �pa��v����h��b}[���s�	�����@�v[ڶ���~�[�wE����NMfV��VǡCtk�}W��ѻ�e���d��o����仸7i�~a�,_לY�"����!�욙n�͍��I�QS��Z�cd'þŵ�}�S�/� }D#�sn�@��"�4;`��:�#CD��?��x�	���X�A��Ts�H�s�?���(TG΀�D>uD����������|5Yv#�G(ȽF�:Ŝ2��w�Fn[r}�;��{V�c�E�mr������Q⫨�l��l���X��t�*�.s4e=��p�96K/���9��uu$�SW����yDMdSzfS��Q$���+�+ޛ�o�5�"��`�
�W����N��Ƨ���$>�s �@��]h��FR(�����	٭�$>��!4codi~�8����ɦ��%m�?�-cZ������� @R�9�i	�8��t�}�H���ÑGe �h���QX(�=Bc�T	9�8|��Ab�޽>�
:l~��Qڭ���|���1�.5W]�Kα�q�b���7��ט3���ѱ@��T�l�e+4X��3�ۂ �m4 ظ��^T��A2��11ha1���c�ߧi�G��%,�(�fs��fc��Fa-��n��l�\���#������g4� *c4����ff9ҞIa%��?��Re|R�-'�#m>���B7Y���7=����GɛX;�3�}�3��+1p�JL�+C �/����?x�2�>q�:���)G�i;y �8X,�:*;·�k�{_�޽����ܰ�V�xW4�:�����,U�H����	���J�8���^����o���*�aڒ/�/��&盢�YS�~Y$��ZM���a[p�@�G�nk�²�`��D��P�?T܌�3љÜ������֖���,�G�Y�F����7��T���A��Ϗ��CM�"]I�H��m���]g��G��ڵw������u����Ğ�Z�h����n��Ǐ��`hW�hh�(\q����b���C*'��B�ۂ�}5G}�I�.Lʯa1�ѕ(B3�ӳ��kxS�ջlZ,ߒ���mVԕk@���@�gZ���F7�Kí��B�12�Y��)Z.���Z��d$���	fvzʟ*�[���	�-�o�8P&o�y�.@ۃ-�Җ�b��j 5�D��-�8�?k��]���Ѿ�ӃΚB���he������h0B3�Q���+W�d^�^!Υ�O�\�˽�=���)f���b���]t��\5�>��C�{��"����#F�<��_��.�ٌ�����Z��А�b!!�U�N�>kЛ��9G�@�PX�	������/��S��Ϧ2\ꃎ�n�
�b�?;.F���;P��9��ӻ�������~4���x'�;WRk֙��*#|(n���M����1I��f}�V�|_�`>��d�e0%�_�Fw���h�,y���J2�uj��V��IvWN�e$��l�p.n���`�3������*�h�5����gU��V�"� 
�5��ѣ��\,�W�J�\����(�<�5TĤ�xF�^�,���
;�yi}1�O�4�EU-N��?�.����Ou�_ł��9m}����tU�b��;�|k��wD��f:p��jc�3	�;j����t��]� 8���~D�us"(xnH �|�L���E=7����E=_�eΖ���!4E���mi���n�vƠH'�
oDh����0��L�VV0D�Q��4-�K��n��j��=85���U��j%=���\N.�r5|���F|�Os-[h��U�@(�X+�hLU1˓F�f�z��tPM��gN����RTޑ���lCr�醧���9"��Ә~zC���M휃��r��vf����<���ă�'`Rb)*���<�풊#���g�t�}�鶵;�����tM�*`�1w��(nI�n���[0z��o4&[լ��/��p>��a�?��Zh2��^(��#�a
���\���]NTKW�2����<V�������~�ﱬ^+㚚���v��%���m랄2G�K�snĽ�QƏ�}�x7#��B2?�7z宴
8N:GJ�G�ȁ�R+�4���/��뤻��!�Sƕ` ��\痋B��k�z��Ţ�2Qdäa�e����$ פ_����K��4@�����+�  Q�N�Rs��0�C�[٫��N;���;1��b�LL��s"w��1�߬�<����L(�휽"7�X����(��'۫�L��#�%�f���6x���1�}�������d5�� :f
r�5C]^��[����kϩH����0**�^b9����ɺ8�q�p����Oh{��6�\T?�ULvg��ѫngn^�)y��7,�h��6[�X��t��^d�'w;��0T�*��R�>��a^)�].�ez5������>�3�f�1�Y�9K��@?D�xD�i�>�����N���.�4���&	UD|��S^�2r��%#�ј_̳������P�S�Y�"62��0I��dռn�n��tb���X9��x��p�ɖh��-��u����,b�o&M�k^�g=�tp�"ۘ �(����Uޫ��g1Xiw���V���E��!�U"���f�8)gƼV���f��'�r��絖5���İo.��'�u�rL��xR7���}�i�l��9Ϛeؖ[
 B_Z��r�豰�i U����h��KB�X!H�P9��Mi�X��`~M/���R*~ҫ��?8,Y�Kե�!��ZP����7�41�|��r�=꘎X���<GŌ�e��0
X�,G֮ox�a_��.�D�bb�g~���םs�����W0�䳜�m:XiN3�\(�	�|�>vݡ�KN��������IjH{���r�<`ݟ�$U!�3����I�E�n���^S^����C�c�����yN5��:L��Ξ���.���׿s��ݞ�#n���!��)#|�.*|r1�9ڦo�ܵ����T��1�hp�3�a��=&~T��ԒTuL�8g���.��o�к�=V�n�Y�q������J��(���6":3��@=��g`͖f����Y�����bcI�]�l2[��s�ud�b�A?���_��{3i�ޅ�\0�	6}|絫xP�R�BϽh��F��PA��0��D�j��]���M�)�9!O���}�k�ڌ�O��w�?�@٣ʫ�c#Q�T������ @���g�����Q��&��x����?�LC��;w��t<�V�a9��4cֺ���8ł��Ou�!(�[l@��Y��n�WZ���J����z����uX��Ը#Zz�Db�h�zRHK� �ˤSP�3�Y9��|s�,��X�~�ڋ��Œ�]�bM.;�ȑ�[Z��b��(d��02qC;#�2 ? �C�(�$�ºdͫ��A+|�ʾ��
��{�M\Մ�&G-C�V�(�Խ��lC�jw���OJ٢�:iE�i��7S�w7���(bet#	X�\�4��{2<�7����wΧ��Q.]��/̻�>B�^˂w�w۽Nc�Zu+�l��D���N'�x��B����`���@��\N3�0'Ь��|���a-������cWLY�[΄'��6��")d��z�p)����]�'�_��<0�u(�Ĉ�?y}�;4D^q�H��Մ���DT�Z������b��[f�"!0�ߏsXkq�GA�`�uo�S%�����a�ۄ�z&���i�i� vC�<��Z�M'�~�YϐO���� X�:md��YX"���I�&yO_�=AP#KO�!/N�����W���݂�㏪��#?�,�vỶ~��O_����V@�d���6��7�X�
����`�t�٘a�_2kG����V�/W4<~���lg@�[5m����ʊ,S��3@�O�rG���"%ɡ���9�c�gB��p���(�%�)�d��3�]I����?F���;�󹾪�H�����Ԛ+�ϥ�v��D�����T��]Z��$=�T�Ѭ>�ǉ�ΦNv}��(��,�ZD�D`�j�a���j� �i<��.�9�*rD���er�	;���?�u
p�Dj�<cP@#�7�� ���7�Vyz8*�����!ul�O��\����	woI2����KG����~+�T�٫/Iy0���kN:���7a�����B��yV(YjJu���N' ��񨔉cq�[RR7{v.��v���h�OutU��Tw��sr���%[��<�3JuF�7�t�X 2KY='��VI�,`9���|�v]��� a"��Ac��Xr�y�!V^��0C_ǆ5���A)���p��Nw�(���T���;��(�̓�I�.<�����&�#@H�6�>2	VV�R,�Uؾ��V*_d��L�bvV��{N	��e �H�2��g����dS�~�e�͈fP�O?p'ܵ��!� r����&8�J��!O��+w���:�-�t� 6��_}�K~�³��r��k���2jMǬ�fW����׈;>�ۦ�h"��\ Й���x	����`��w���g�z�He�
C��iui*O5k�ѸD1��$��y |�aK�����	��꣰�t9Y����b�_����gl�G�vn�3?��B�0��*�"�>9/��	�E
��)�[�P����T��������A�<tC9���g�Q�zR������n"�J�j�H�z�ݰ �<X�����{7Oާ�QX-c�� V¸`�H/�E�8���&5�f����X���k���.��3��>�w��6����-F�6�  _}��E��LK��C�'��6Xh�o�]�X�Y"�|$�E����U�APQ�{H	���v�5����U����q2�I�EB��K?���U�x��|�PW�t��2���\�6¨�;s��+?�7�� 4[����v=��Fc��M����1`3�PqM�v�9�������
��|�McH:������-P[�vw�l� L|��`�V�1�LZ[�6���
�3��i��qR���&XSzr?N�bbzWx����ᛙ^��n�Y=k����,>ңJ��������ڵ�]��O"X�F�(9��0�/>��e�b��v�C+����Y���|�^~�1DL]�qAU��G�6-�~�XO�`[����m3�^pxO���Ž�Gz!<p{#��.ՠ���Àn������x+ኜ��"o���hh�g��Ӝ:�8��t�d���$�>�����&���T���@������e�<�jԎ��0�!:o���V��N#�&���2�t��]�ɦn1�����O�D��u��={�˲CƠ�O'y��y3��R��)A�?`�ڹ�g�1��C�ʲ�DXe��x��J@��	�|z7j����y-��A�u؂O�W��@U��ů���I7H�[C���\z����ve���0!75~�:�!��u�[���I&���7����X�����cCw�`X����Kx��[pC��"wʆ�!7���W��N\ ��l�{>M��O��!
�1ו�=Q?�s��K㝖|@��V�mv��4�*�b��@����;����w$�k���j��z~S!����$V@PS�À_���l'��5&�/��0!�D ��O<�]>"1t�6����z���+��J��hh<@��T�<��号����a8�8��K�ȩ�3���b�>9T�NUP�	"��/;�_��qI�sY`����J B�6�Y�7%�:�l:�+�8'N�(�`j�vd�܃��{�ɴz�A��}.i��~(�?�����ʐM�+5bB�_��b^���VD�!�%�!��qM������ؖ�|1䞂1}(�W�? ���,y��JZwt�8� �,�CŰ�c*|8W]��h�]M��Z^0��"�}GA-����֮��ߵ�~�����)B`GG�}iф����#)��,�34d[�� b{w�S�A�&P҇�T�+0{p����_xQ�aC>�ka��GZ���$�]�x�S�9��C��f ��Wi�T��HJ!&�����a��-ѐѤ���[��ՂB���/�Y����W�}^�d���` �·r�͎�w����1�1�;�7W�6(�uhl1*�0E��k����X8�?�����yQ� �cR�L�o��߶��;�@��fϒ�墜�f^����TI���X*_o��S��ߌ�Nު�l����
@��%�N�*�Z�!�z���LQ��o�B;�0�.@߾����:�.��Y2g�~����G{T��o1���I���'���1�x�l���!���{\�Yu!�JV;�8��0���)X�{~X���0�1w!�.�>k�̬H�p	�����K�T�L2�{I>f�C���mp������h��>-u�Eї"B,1_�C^*e����w^����)�p'�wI�Ģ���ؔ�?ýR��1��J���ÞM�Cs���0:8ah�����_�~\���pO�T�=
8�ة���-CM(E���q�2@�Kz %��v�u�?�Ӎ��	#��i0�l�A �ΞE.�<�1�E��i])l��?61�2��b��D��fr����-9M�>ms�gO�$�K.�UYHNG��!t|-�/���џ����5��~���¸vv��w�;�Pb�V%7�|���Kn��mu�:x���s��ެ��ӭ�*{��agƅ�<��$�L֛O�z>!��2��hFQ^��ߘR��E*����$�����F�Ho,�`����0/S�c^��^����v(jpp����qE5�i/��_��ۚ}m��vͼ�cIq�=*��~M����g��a����b�,��P�p�{k�&۫-0�4���j�7�X����ޮ�m�YoL����v���>�h[F�k�r�f9�,=�pԉ�/ �w[�B$�@�8��e�(���f� =���˽˯��Jf��W��dg��i1aUԜ>)g�3d �Q�j��#m/�ӈhg���F��v|�%��W�)�>6@Hԭ>V$�UU-�j�Ǵ�i"��2�������!kN����Y�c�v�#�p�����|�E��i���>�b?V2�����8��jP�	,'Cz����t��6��j��=\�{�5�#4�w�#��R]��b��@:ea�Pq�Z_�A[����o�����z���U_�B�DU��B�3n��ÿ�|�x�'�����_�̟Os�G�Lw�H�G�-J�����Ac
��aN-6�֜�&V�,ZWǿN�f��pO�Jh����~O��D���KK��3A�����gQU]n{��w�mJ��X����<�b�p$»��[gGy�zk���?D�t�_�u�nxc�Hͧ? e<�Z^��p����%f�`��S|��T�9�F�$q�[��{@Y�N~���YHh�r�{���&�kW�u�,s�ϴ���+�'W/!�����94����"Z�y�QO�W��f�=Mv�IG��u���p�z�v.�.�#��l-��
8�g`A]����}�&f9u�q��b�����U��;���� fw��f�J<���Nf����V~�"�ΨrB��C�i���"���e`F��jD+c�f?Ɂ���
�BD�k}q�-aX�o_�&!-D!?�������2��2��w�n��fw�j~N{j5��ҟ]�S����Ŏ��X�,�,��驣�r�+�ڬX������$T2��<���,��Fi�^��κF�����@����<��v��a�cT���mM������^ʯ��7!Q�;X�.M�U2���M�����09�E��%��>Pj�4D�0t1O�Q�Xc�����(8J���8�o�������j5��@_�����KWX纁K<w�|���i_җ�Vf�ȕs�\��k�����`���C��������j�t�Ɨ>[���`񁄌��vd�\iS ��"�:�P���\�\�­1�'վw.���QAMW��OOB�O<�E
rTx~���d��"�6!O+��"����Q!�f�P��r]�U)�z�`0c@����{���Rn��蜮�����I.T��Ͽ1�wĉ��V&�>��������c��b�cˣQ*�.��m������_���E�ɕ�-��6]I�q��_�5��hh��=���g��y���_�;r_���&����Z�J��H�7}JW�(���dph�5c��+�"Bls��_�m���7��@uN� ��X��Ř�;_�)@A�����&�V�)�ժG��1'�<j��E�{US�o�5���'����� �q�b�/�x(���6~d	�۱}�1b�|���U�C��Q�C%QI,4��8󧚏ڗ0k�Z�p�$��1�U���С��bOt�p�}�3&@#O*�U`�vy��u�nI�Z���Ԃ1Y��kq�xId���m�ȣ�K�7���}��ʐ��¿��D�8_����W,��VR$�#��8��~+��rj#D�� ?�;�*�E���S@�|����,����3���-'���˽^̠(��W�:�R�b(�ke�ƈ�|F�g�\��^�S���u�k���㡫:�]��z؅��!���B����у@=�4\�2���J�����~(*h�(c���o �܂6l��(�K'��ho�4����Qq/�DM��>V#' J:+W*�ֳ\�q��� 
�v0bB� |t�mg����8�KՌo?���+�q���h��xc��H�\��"���]�I����[g��X�ߟ�����E%�T�,�T&O�츚��1��6?�vcY���O-g�W�p�����LY��(4�'ed�E��@%���V��n2�A��	��@y�\�+7���մ�T���Owqw�2�u1����:�Ft
�T�7b�N9����5�e�j�e}��j��,#`�N���E�ni�+�ɺS�l�*�%v��Y�+�l�N��ā���V�Lk�aĸc������{-o���v�p�j=��7˲<`_q6��`�M�6j� ���3��@swn�|dK���#q�:b�p�S�����|�(��4>�7���.���ڙ��N<��&�88��~ܹ� SX��v`γ�a����>�*����^J�.����k�N�_��l�j��u���˯�uMl�=�_j z�*٤G�71pH:���R..��c��q�ב�t������u�1|���Y'\��f1���	���pݖ���Ȣ^�Sa^C��WՂy	�v rރ���0y���Rn3m�lm(����������%��m﹋����A��`��?�/\'��Z�`�>�Z�g�j�1�qv������o�؊hW��n�!��Լۄ9&y�;1D	�OV�.��|�]��6�T��jGq��(j���\��I0��:��'�Yr��/�ev�$b�<�g>`�xb2O�l�V��'v�|h5���������>u�/JR�K���<��f��[�2��~�4���eE�?נ�ݮẂߤ�7=���k1�)l)Q�4I�'�~������66��t�E5D�?>�.j�݉A��t�N@N��:i 0U�{F��q���楤`A��{E�ϟ����6`A_?��G���Q��cx�8s&?,`����| s�madU�+ڬ�*x�o&�S,)q��������Z�ۙwԠ9��JX��og�4�,Y�q�v�)��c�.ko-s��Xj��	��F|�UP�t��^jv�q�A4��!*��f�ϱ��F��'�#�m��?��W���ۈ}�� B<c�\�5щ�OVx��y`$�5#+�@�-*��/�R���I>�9�_%���]�恛����W�:�γ�k�EB���u����.�pa<̥��)���w�ߴ!�`�����ڿ��G�O� C���k�y���n"k>n�Yo6�����PFuY.g狣D*:v�pC����z�oי�\�����8mª�
�؎ �� Уv-$��0�-�;w%��`R7���S�4�ӏ�.�^m�i,	z�!9�o���}=ɷF��I�9��ٰIMR�&���Va�M�غ[�%�Y���+�*Q�+s`MaK����I��[z"{�k�u��o�T���!��1Z��$���ܡ������@�C�Cs���LQ+�2[�����+J�������]�$�7茲��%�����x�ŗ�A-*�^�xp����,�~�v���aׇ��#9 ��D��2�J�?'�E��ZV��-^a��as�܇iH��m$'��w�[`���0��3r��ѝ�/[x��
�%޳�]1��2@Ok꧹DU8?�~ى<S��Sq�O�nפ&|(R��D<*r78�y�����I��+���>��&Vϧv�ܺP�����x�yס<���71<��߆c��Z�}3PR���2����s����z7�J��8��,d�nH�*~��uf΋�f
��x�!����O~q�al?�_D���RZ.4)�f7#ŧ"A*iW[/۴�Bz�|�h2�w��.5�������N�EF�΢̘�1=+"eP�h�#�X7�)�E��H
DJlp �8FJ�N���C�?\$�1�q#��>��뛳��}�HK���g��S�h���,��շ�!D�>��d�qԡ'
E��a�N���H�vm�gb؊HW��Gʶ�+{ީa�z�b���-���ے���A��D�OphE���T�D^#'�aYyK��0���L�ג!)��N���@�[KYm^3x�N+�� �>������O���U"�ה/ɓN��}��fX�{6�\�þ����]��qb5�LwIޘ����p�V��d�_�J��}�p��q�h���?�
������z���!UE5`���ڽ�I�1f=���G��G󆃛�=#��Ӷ.���9IļVӛyA�%�~���#�`��s�q�_���A�NHCӘ�j+���PL��G.j��i�����e�a{_������yo<�4��0.����Em��G�,Q2�*���)䓸�)��/���0n��E{�"�녍�c/�+*[�&�����J�L�,�ɪn�L�}gv�劄)�m��1|���?�3�pDW� ��y~��SD+�]������dT�u���n�ڋ%\��Ѫ�����Ĥ�[�=z'~A�⁣��e��Tӽi]�d%'ʿk��=�IT�r��g~67�?��h�^_6���:�/}�d�q���5�����;5�o�-D	�p����;�B8��O��H������xۃ]�2bK�X�������������jKI\���Oq��q��K��f��\�$)�����c+i3����;��̻��-y�-Q����K���[�q$�TU�*�?f��xR8s���扗lp�L��r���ڬGل��q�H`���"��Et�O�ܗ����$�D'�~�NFh.�:ЎN�A��'�#cC����Bg^��m�1�U�U;J��כeB,�p��M��~%�ON�o&ޘ(x��<D\8CM>l�ƿ��b=����^�t�-(��;vǸ4�*Q��Wh�"��9�'9
8�SaG�V�æ2Ձ�UI��C��8M9�Y;d|Q���
ժ˦���fQ���`��RKᶋ� l�t�`\���)&�m5�8��<A�Cu �SԄ����&+!xi���m��4�q��3�iPJ��hXiPy��fߔT�����]{ڕ�.�����u6��w��u�&������^���y�d�����y���-)�=�}�͔�|�!c���e�������`��O爸�{d�Ե����-��;b��1��񊂪��`�EĲ�9��]ƀmԌ��	�%nL�����2��]k*��8X����j�ǒ �Z	���P�qA֫���hv�V?"��m���&�\փ�W��;uZk^��٣xқg��h���j8�`����f<xE�,���T�0c�^��@��?��\�L�S��W�lާ�N|!3Il�T)r��M��`�x�&�`R˛�����*����rV��ՠf]�ٕ��!�j'!<��U�o�}�d�8��ޘ��[����e���p�Px���и|ϧY�����9�m} �1��)X@��bĦ��+g��U9EY��y��hz���0��FK~�?�L�舗и��@b����j�b`E��rA6�2(�}��UnO$-�հ���f*P;0��U�#,.H��bZ�i�4~��~dm���%F������ddՉ�R�-�<`�%\W���������x�I�EA��l�'�{�:�?�e>�Af %�q�f�Z>[�g�W��,�lŞ������&�6���̿_��D*y'K�d�)�7�Y?�m�j�I��&�,;9���gWyF&�f�/D���@�F� ��ت�<���n� 䇣-�������9<������0JQ�O
��t�I��.O���W�^n)��ߛA�6W;L�sWp���'=&y���A7rYf�d傔����}��ͰXsFQ��V�D�8��3ׄ�\�ګu��xG@ʇ��n���$D�U�C��C���G��3T����v��3��̲�P=��� �J�{���_ ;_��f�HФb^��捱"Ҧ^���̬�.qP|���v��EO�����Flܥe�S���h�*-��s�/���j� ���䖏z����z���ר{)�S�s۰�(d�8L�?�O嫼��W[��x��������y8�W�"���uϣ�n�ֻ��Y9�H�kH�Z_����G�0aK�����-��y32��0<�f���33�l��愲�:
�b��@Ul6P�9'|�?W�Od�	<��52�.YbQ��Hg��վ#ZcP����<3�0�}�o;�R�"�H���5}O���Uݭ���"�(.K.����&.3�@��<��ۑ�TQ=yx���(o�~%�!���l�OX�L�'�K2T��0����	@���^��;8��iu�W�����BlC̩�l����*�������b��Oe��x�<�c�P���Ū(@>č9m>*����ܢ�l��X$�exw1�⮋W�����'��:�dި �X��!��Ę���i;(c@�-0��/�̝�1n�r�?5�W�Q"�����fL�O~����y��A��9.�XG���Mz iV�	w���/�ϧ���WZ*�P@Z(���.G�HBZ�I-���������*2�ċ����Re|�]������9�Hݏ�c���¿��J0u�Pb����?���^�kD����k�'0F2r��O�3vi�+Vi�,z��,��:�(wdQ�3�Z|ٛҽ�؎"S�e�ɋ����6���"2?���-�y��%@���pR�����݇& x��o��k��*oo��ӆ@B���{^Ϧ/�C� �:�mMC��1�"���S��Rܯ6��1�)��"���F����l읮�E�%M{��fv�8�YQ^
�x�R�~�a%��LO��}��@NW��T����iU��>�j�b
G��Ǖ�M8�c�`�VoA	�b39#�v��K@� ����;qg�B��P�d���]uY�����vl*t5�H��1�}��3�^��j�~�T���k��CQkڌa�w��4	����	T0��rpA����co��O�f��e?��uS8�P`����3$`C����:*�z�-���j��l�m-���in�����m��4o)�)4:Y�'�8��_P�h�t0�6��/F47��I�r����o��	�j~���z�
*(E7����*"��b�n�Q��E����z�=��sb)=��	�	��ݰ�N�ɔ���Bm� �6Q��W:�s��z��2!|]�G��"#��*-U��Zu�L�2��f^'K챉��y��(Mɚ"���o|�6���W���(>W��H�z���PGr`��J�',���#I�`<ǣ�};�Y�WZ0�Q�s�? ��h�m#�ו]U'ц_o��1u����ٽx�P�8� C�j:���hD����t�o��i�5�*q0g>7�Ge�"�����c�9\�0V@��(
m�O��@˃W�F�}j�ӬF���Q�rh��B�6.0�����mA�2�R��m�ރG[t^�Ω+@yd��,e�q�8��ĥ>�շ�\�[��O>�����>
ö�:��(>,_�ͮvΎ9.�<�4����W��~�P}�S����e`�A�W��Qp  �?]��6����O�C[0z��t@�r�I���J'o$b� ���@�'D�	1���XNY�iߴC�*2��wێQS�DR���0	 �8��%^�P�4zǸױ��xU^�?�l�6�=�f9�����-�DeM�@�2���r�Y'�l�gK�M����2:[�O  �����O3_�9�:�da�,.��1���3�ޗo�l۱eDC <p�:I�N���"xa�`Y�]�"T��?��/�/B�~9��T)�J�ͻ�Ɋ��`��l@�i��X���5�H�4� RZ`X�F֍��d��>�G��n*����8-�~�>Ff�̅ױd�g�ɍGreƢ�x],v"��`�=��ĨJ
����O�(@@��Ϝ����g�n��(@�N�����?I�����>�^�w^lm��r�9h �2w�{C�q���6�@̈́&��z��@SI���W�TH�Fxy5��`9��р�ûq�{i�|n`H��#��p����G�ow���*<A�YJ��k��e<E��٪��t�ǂ���G�ie���G�����50���ñCx�~��Dtu�O�Lv+'4�yt�<-}�f$��%Y�*Rkʾ[B�>��wc%AG��K�_3�G�ص*���g��GUY�Y"3X#8{hl��r{4u��3�5�0T���|�	�-Ccv�ɀ�$�|s(�[��*�Xd�Cf銻=�^���|��}Z	:a)v}B!%��jqF��=[�e����oS��°�il��D�?���yK�5a�_r�;���CL�g�*��1���\z���/J!}t��9խy�f@_�Wb։��
�$�OCz�S��
��L�R*-�g]�'��Wq'�̺�A�� �ׁ�ZfQ{LmE���3�2[�S�K��q�<t������AȬ=�z��hl������Q� �l�~F�UA|($�/p:���N-Ef.��ȋ�%�y��n���~�ퟮ]|��Q|��V�	"���z(2wf�X2/��D�	A|���1�s$�j��o{V�'�*�g^JE��ϼ�4f}�cM�zcy� �hA��⒵|�g(3��0� Oe�q�Cްݘ�xCҮM�����.?_�76�j���ⰍISs3��X�����o#x&ϊP*D�s�P$�&�f!�E�1=����U�=��Ω�Px�k�sq[10`��&$Ă�ٵO*�Yj(���\m	$�"��1�O�������RC�n�	��n�v�p����'*~n���5Ln��g�n�H�d���99Ԇ�.B�ն�� �:��C`k"�h*uom"����UuP�kIS�x����Ms��O�U	W�X�P ����E���o�H�A�kozxI�������W��B�\~Q<���}q f�ь�����5u����gz�.�$��M�*Q�Ϙ�����K���3G��|�R+�B�4Η
@J'pʹ1|�e�&nR�^U�aȕn|����ß�D貊\@3�n�ΐ�\��@�����S����|t5	8Y�Z!�8[��J�fu�-փ8�-S���-���C��èQn�O��V��L&<���A�:E{��}h'Xu3ۊ�ϗ� �f	���7�K�@َ%V�鐉_�	��O�[��\�^��k��K+�_Y�#��e���l�v �hޅ)t�;s(���tH��~���<�W�l�?��dݨ��`���8�����
��'�q��.kh ��S�*a� �����6r�܂ا@JvB���@�?�
,�w��D�G$V�zXn��UX?���o�{D�C:�;�*Ou��1�8}��A	��6����{��׮�=rd�(��|��P��@�$�[Q�Ñ ���x�L ��G#� �4\N����7�E*|�uT��S���Cs��}��^���e��k� �dI�K	�V�_�IEH&���%dl�O���W��H��#~f~8.��-O��8�&I��}3b�kL�. �=�(;_h�M�t1k�
,K"�%M���l)����DF6��.�#�]�n]��K��Uq��['��
G�4�������#P�����k��G��4��fXwc8l�4�-*�I~���:�CDj��N�^����$O�t����I��:�GH/y��v���1A�S���Q"-�VP-*k�d�!�E��&��òc=���攚�:
Rl�nll%ՊcW�Ĉ��pG�Q�-��#�����!y�s;����oA��I����V�pͼ=`��k*�W��lx��t�Ǎ@7�s�ʷ���b��P��1����O���`-���s�e@����� �5ܺ��|���z��Y�+�v�2^���泇�'p�HƯ=~D+��:�P��*	+p�iN츹�h�½P�C5J���n'bMib��a�4!p��x�m0�&&��3� Z+E��%4�����ŁW�r�[)+w��A6)IE���s�rq��>L�˔"��0 ھ�F!�ޗ���y�໤���Ժe�UbÊ�#�܃�ʤ�O6,'v�{�R�1F��M��j�{P�SD
�oE-��Qf)��%j�Y{�@��ƒ����N������o)l�9s�|5qB\"n�]>L)_���#dӰ֥}��5�f
@��˽Y n|F E�|ȴ���@;���#��n�k�cY�H2D�COe؈�j�ߡ��т�����J�&� �@����Ȩ_X]��dV����W8$$d��q���fR�g(5_�]���?$�9�G��'Y�`�223q��L� �|��w����z��ᏡہwM�&<tV4"f�h�Jb�1G!ܸ���uu��L�AU��m{����������bɟ���c8�Ŵ(m|Bŷ�;�I�Ȝ��B�#+/�(Q�\����x�X�d͡��'�N��I&�ף3�M�BL��Pqy%��a���g�fP���ԉɞ���c�����7?�)sJc�8 �TZ,I�-��K&p�(_s&$��`�$��5��{8�m�M�[���m�i.w+�>߲�t��7�<��"��jFĖk�����,3��Uv2ݿ=�������e�I�t�U'�l���m�r��p֣��m�ͽV�Vw�.���t��]��=�Ȭ��L�E{��p�|$�w�k.�{��I��C�����k�OI�}�qh��?�^��r��
���P���XBwHx��F�����̽Rw�n��?,�h]���Ce���}]H��jH#��n^E.��d�[8���k�ه�� �Ӫ�bB�
.e�u��P���yW曼��-�yfz����geÓKH��'�u$���hh��w�nbN[%0r� ��j|a��07�=sB�C�#�5N.��e{��|A;qH>��i��/�n���V#hQ���^���Y@nc�h�n���Ky�ϩ5ϖ-����주�30�6>�:��"���$���!W�U@ʅ��lYn�m�g��i�uQ]hL�(�3}ue0�|�#�3���B�}KS�������'c�©x�n}��݅����z�xu����ȹ�m���������|r��֯�R���!�T}�����ld?qʺ�ξ�c��B#��nh��o�h��O4���&����jF�2＠A�5*i:�1�Jx:OQ���D ;����(	Fl�Ab��;M�B�ޡ6'��i�9G�Z���z��tq���!�����u�ު�c,-BM��q��.�#����Єp� ���(E;zH6p��z�n�Rb�Nְ,7%���tL�Fk����M��A^Ŧ3�rn�'���M�G-Iێ�#g\��.��ڹ�9߸�����p��q��ѳ��,��ի�@=j�[����fs;z�8%#l����K�w,A��.��ޭ�O��b_�H�׻�F+Ӏ&��1�/����������L��r�����+���?���u��k�*�M�l�i#<��d%>���6��v1�z4�V���N�T�w��L�To���F�`0U:�|3�(�O=��%�<�ҞhĠ�V@<�A�H���dy��0C~��S^!5��Z܋����@�[$x��*�7"+�ꫝ�F�4�Ɔ%���	�u��eB�\��_]�c���4�[��pi���m���V�̆oڗ-%�w��Ym��<�XG�s�i�`S(S�50���nC��n��R�Q2����b|r�Z�7�Q�UQԮ�U`:��yف��M���$c�*Ʌ�#g"�2|����!��C���5�;�A��ϲI�8:y��[���(�J�nu�ɘoL� Y�Z~~4�xqb��5�3;b)oZ5��ԧ{K�bۙ��@�g������W.o�ɟ ����%!@F���h�E�ګK����k����"�`��t�ȓ���0�{B(ͣ�Jr>�R�@�á��0wi��6��m�2N6�䛜�j�t���N���/��s���r�,<���n�mT��X䢛�U��'���|m�`ܚ*Ӳ��]�ؕ�m������|É/G�~�#,���r�aaxpWg�Nv@1�V�.�ꪘlU$�i_P��#�^(u��P���z_p��܌�����`C4�ֻ4#�����;��.�m�Dt3��&�%�ŉ��� ������Sߣn�*�Wr�425�hp��U�GUsb��T ��+���9K�úPC=)CFv0�OX6#��N�P%s����(�Q~8Uds��`�졜�6zPF�����D9 ��=��h�'d��X�ҾD��(V5�pD�Jhqczƙ�e��O�q>�(��KS����pc��H���'��5�����j�b	9z���J{�	&�AEW兌�����៻��u}�	;�<Qp�&S�AK䅃z3�+����O{A#q��Xm��n��Wt��HW�X�	kE҅�m�+�����|��I�M�)4h�}�vcJ3��8��T���+8>GM�[.�	7��]ꟈlB2��iڷ}��Bfם��b��WIF+�b�56Ɖ�2�[��1V��|�_[���-��Be�U���(���`Hk�Ηyq�^�H�uC4<����źو��|&!,��	�s��	3K�͝�]�u�͢ɏ@4�k�e� 05�d���S5z	-7��F}�)�8�b��2�n����cƷ|�P�!�Rd��:"(��U��S���$+�� ���m����+l�m0ȨÝ	�)ݗ�)�T�>�2��r���\[E*���ս��Ǜ�>�����c�!��$�)�P��"��q�E'���F\�W\~���Km�#?���(d���I�Ey[��)��wm�<P�� �LM���?H�o�Q�����r8j����2A`��V������E�CG�n�DD.< _���� M�'��yt�],Q^䱧�v���'%E�1Yk���BȮP,�p[�gg�$h��@�rI	#5���+Mݻm��}>����<�uQ��}U�I��r� &v���-1Mei�cn��C�����*#�?C�.�/GR�s** b��������y=u�L����v)M�`� ��d�/bQ�L��Ŝ
�A�f=���������j���:��9;���_�4���̪���+]�+�r��Hp������&�9L(bHh�����ֵ(������[����k��a�aF=��l�Q�bPs�4�~n���/g���[�O=H�C�$���P%]ϳe�������	9а���SBR�kV��Ѹ�n�yp�_��C-�uzV��q�j=��;�C{�L�|,�M׮�U���TS�0k%X��z!g��c��P�f��d䲥���L�\׭�Ysi���V?�RAK�,�j}�\c΀+rT��s��3�a*�:�;��"?�0�]`�5G��^,@"ƴ�ےFi��S���6n��sR�_��H�%_��`K聘L'Rhؓ�}�^鲢oX$�\j`f��0�VԆ�4�/�Q]~g����J]�g������p+U�Z��11���=l~���!CO�v����@�*���Q���BC+��MQ]���J�R�3�<�W�<�qܯ7��c�<�U����E��<, ��o���F*�o�!���Y�Vx��\����X�����-q���+������W׉>.���oW��:>J����_]�T�y���OQؚ ���Q��u,��7��;l�L;><�+;>�0^|K4D?�L5	�U�"������?�ٍ������OP4���vB_9��V��X�M�n���dGp���n�m��jls�-3�J�o����D�fM� )r�Q�QN� ��Yh��w��̩h��RȮM�U�k�+�����U	2����w�l��%_xD9��e��᦭��fn9[�pdR=��_ �N����^��y�F��Tl�Lb":�k�Hkt�� #[��ȧ�Б�i��=ӥ_�ij��<O�h��#L8�*�e��.�!!� ��oJ;X��i+M�p���� �����7`�`I�5���%�\�d�ar��>��8!�G (2�s�5[x��0�vtƷ�7���e��bM��9e2�M�.<Q�Ѿ�/;�R����v�����KD���)�Y��;q�k�<CC��I�h��
���4-�-��Hi-�*� ����zW�h�̪�h��d�<vj{��%��5�e�d�
E�G�޵����Rgc�Un��)��D���I���XO��`na��6X��Ҕ#f3�{0Êc����I��nf�;���NZr�����wXy���4,0>oh2��08Y����~��$(��� ݨ�f�׌J;֫4��[:��GE��޿�ꅺ�m[T���2��E}T���o,�Z*�jS��E�4V1HCߧ�X
�=궥l���繻C�p\�Ul�is{�6	��jm�WA�� �j�+j��>b�rp�N�V;���,T!�Q�$ �}eq�$,�������P*��|a��p�*�TﳓT�%�v���>%��)��w~�[���W�:������Z^������G��9<SacfǺ𓿒Lwz �7f=�9^G-=���f'�
��o:sx�������S �X�C_�o%�}���	9��j.C��H����7��%��=��gu��S��b�� 8���<�'jA�o\K��{]����(ݕ�[��g�:���1�1�yĝ8`��;�?�k�Ap�.��9����p��O_B5��*�$;$f6B<i��'�U�XV����U��|������@A��~��T�q�/��/P�+gPό�)�-8�(o�֖Ś���3%��Vkǚ���t�����
hǺ�a�bр?U��g����Lru����T����Y���;��iͺ,��/C�=lT���d
��a#�z|h��MA-Jz
�S�h�M����}�ɪ�|�&�w S3ZlgK)J�����f+�4�	F��;;`5.\����~̀P����;����f3�.C"�ƽ�@�?�T����Z��@��AeKS���@ƠM���F�5��3ث�2��GްS�&
8����u�'�3k�sZ��ף/�̟���cMAR|(���p���1�IZ��<ubL��� �-�8	��_�VeY����B�v�ڠ�#Ć�\2SkM^�y��.9,�ZT)�,�&��۬mi
�0���=S�`������ ��N�,ɭUO�=*Do��0䘡�h���m�\�|1O]V���0�y��-���"�j�'�M6*ξQz
<ՈvʱX�gP}oADؿ���~�щ�5~�]Em����<f5��ppz��`�}7�n�I�[J��8���7��鬟7����;�V@cd
�%luҬ��g��.u�u>.�� Y�Ч����/�C�?o���Y��	��m)�;Y���e�v�w��@����4�4��������{Ǹ�p������SѿG�&y�"���B��b���ż1�8�|39�ҧ�9��A�R/��U���	��2$ƶU�<�[���,����"3���@�	��12�HKJl� �.�s��"vҷ4TB���һ#D��D���m��b��@��Y�\��j�#���
�f
a��/ť���<.<)lqf�׃��� 3<	��C��(-����gg��y�m�,��������&JQq��5�&��H������61\���/�¦즖dߧ�xm��¦���X��/��ۍ�Om�L���}��usv�EFlt&�d�寧G8P��mM��u18F賽�5^�?[��t�(����8�y���/�^��Ma�j�MR�)�?gh�&~a��f_(����9���l7��X^c��c�I�U�n�J�w<�+>�gS&�����A�+2��aȽBz0]k�d����y�"�q�h�u�����O�E�A�F������&��z���3�&�Ŋb�u�[H��4ط���E*�	@yØ�-�E�R��]�}�&�8���,֕!�L�e�+9����K��Ar�w��(��/�H�7�TD�R�qBtK��x)�g:�K�+%?;�(���P�(�'�R��D�Xѷ-Cѷ�;�/�Cw/��ca���9��&��J(�J&z6�����Z���q9��9Ԑ!�����piG���A�Ҏ��$�̜��'�C�Ȕ�DL%��� �۶�Q�bpT)΢�d�i3��b�3iW�}�U��^�m
I��ĔX��.m,�qi�q�⾃ז-_��Ȝ+��E�!���㆑ǂ�n��x�q1�T�C��EW�~
R�?��R<�pk�Z�fC���H�fކi&�!d�,BF��R��?���iby}� 4�&���ˀ'vT�2�Mwlb.(������>�(`C�0��"6K	���%U��Ȧ�I��|�6����y�~��N���>roުS֍�dQ �3Z@G�'8^?�Zǲ)�J�%H/J��@��ǍjR�|����Y�����bx����z��J�жM$�J`R.������*��L�i
 v��jZRРcG���A-��}U��*�j���Б-��
u�Gr�W����" y�E*�	z�٘O� �)��'�-���2&ā��O?����gy ���2�5B<{�~jd�Pe����o'��f�|e��)g��	�����}�`_���_�F�����ڙ�����j���۝C�/�v7���T��F���=Q-��%�/e�3j������ЙZD��cz���(ȧc0�\�J��- ��R؎��@%��>\ޜ.cb� �q�T���`��Ie�A���Go��L#rkY�V���|�+i��qͦ\OV��$�
�|Oc��[ v�_��O���T��Tpv}�9pLv�"bM�(��h��V�%���*�E�8�ҏmт�yb���=��S�*�;�R�;W��|xcGT\���hꅼR���^�+�p5�zA����d�����yE�SX��������mF�"�z��jq�z�3/�����7ö��	��<1KY����x�|�mq�>�ka������g��w�
���
�WCNcA�s	������ӻ�ڋ6�nf\���Y*��XU*JĜ܁��*/�*��dg/F굕��P.e�����t�t8S<��`��JNSnp%^��]N���G�(pf���<���3]
7��Jʵp��O�L���w 5�(�Ev�䖔 6�r�&�B����4?��z�**��h����)Gg�b��h8�.TۗA�i3�V�Wѥ�b@:�I�R1�XW'�j���Y�X��OĜ�� Pq�˕�q��t߽��&�H Lm�e Uv�#�nP���L;��m/�*��l� Nl�+S��K�˥������+e�.�5����g�M���>N�&A����Y�B;���5��%N]�s	S�Y��@K3)��2�ZE^�U'�ۣz1qF8^yz�刃#$;��!�U�����M�9�CCg����+lO�$(���5��aj0㈚�U��{8	��[�6���(�W|'
�D[�B��.}�5��y�q�9
`ZW�O��[d�Y���1��^AWiU�Y�VG�(݋�'=���k���q� 3�\xD�t;A�ߢ����
�
��6��xo3/�V�'�@��e6�x�D�����tqOA(�(l��r �����'�>�"o��@A�P+��-�S����a�V�[��ni�)���^�r��Ӡ�e�Fu����ح�R֛����t�d��n���$t�E/x����F��>�乷r'o禡4����)"+�[�8SW��o	�}�;�a�f��e�50�1R@���tO�p �K��A��Ǚ�b���i�����0�1tQ���+���-����c�`�.�վ/Φul��*��$(��d�n%gI�w2�����x�B6 ˞��sH���A�^�[�J����SV'?eVx���4Y�'B#��2 �U@^n�͜��I���9���_�j��b�]X�>�e��8���f{����ez�n�S4�<U�5�W��6z�0eN)d~d�Ȗ:f���ԛ����f�ʗYגFF�%�b�Ǻ��˽��97^�	�����&m�6�Hnk�)����������8���^UĄ��T	�x�kC#>�n]�GG��آ"z���*_���.�X���-�������#�L=D�?������V@�'�➡�y�6��h�1�E��Ǚ�.���Y�k{J~:V(e�2[F��򋺚�U�Ǫq}�N�Ͷ7C�g��J��YEv5�����6v,B�v�K\1RK�w$#j�W���sPA��U�n�<�-y�eJpj�����J��;�����0DJ���6���sck=I�Ri��
�ۨ|j�T��ک�0��Ac�A��N�]�]����A�ҏ��b؂=����v��Z�'�]\%�B8,c�{n�d���>p�h��L�T��uF��8e����ȣ�,��z�
X�>�0�G)9U�xt�-�X{R�+r�j��$��=���O|߫`&?"�I�M��c?)G�K�ʨ�a^|yO3{����x�ҙu�ɺ��M<d�Ә�Q���+�o��"�Nm�ղa�VJ��^Ю1�j9n������������*dh1l4/���b@�������$O���DR�ˢE/��AZ4��i��r�7M^�kC�$�*��cn���ɖ�7�+Ϫ���g�0v�j��WM#T(^g5f�=�]Mq�x�3m�R²-^�w�ߠ_�98��1�Qr����]d$
��s0�ݓb�Jh)� �[�Lř#W�jأ�CE�;ȼ�x˔��Խ�{]C�����;��H��8���-�Y��Y��-��HY��F�J��^Y�[����Z^��O*?�平��;Lz��\�G-�,	k�[���>o^�^G�I&�x�������e�`�t,qo+d�X��O�k8m�����
��԰D%����<.�U��rQ��W�؇1v�5��SSt� h@]XQ�`�ѮY_xWV�^�����zs']�g���
�c�Ȋ�8(>�ĵȄ~d��;�� &0�� }7��|�RF;�Գ_���UtB�Η�>m2~�Q}|t�.1���%���\�� oFu��n�@5k�Gq��>"U���'<��1w�V��9s>J<B�^�����m�gؿ&�sE}�vʙT�ы[�(kl/�~��h旼�0�[�3�z���&���n�3�8���8�!��y��N�6��n�(u7�O��-⃴�������Y�1�r&8�z�rN4;�:���,P�L��ujD�*�}�J]�w�,�:��`��|8�R�}@B�H���|�2޻ΖЪ>��Q�*�-ĩ�X��X���r��zm���A&k���<5n6�'�1��$�	�V�t���>A�����uƙ��eӠ�w��E���hL�%���Ǻ�3+B@$W���$�a��R�m ��.P?oa>�r�� ��1y8�אc����3q��v[G��_w"wK�f��ҵ1�w�qPM��\����?R�8OtS5�H�gOG���[ �$��<R�!��FGw���j�F 7��m�L�w�ʙg���l�y���2��r)��۵$�z=�]Q֍�v����z4��F���6�I��1<�a��ڨ�MC ����s�n#^��?�_!HSO\�� %��O2^����m~��ٓO�R�sC{����ص�>]W�����{Cu�A�A!ϻW[ꙞA[b:�+�S`hѱ쳠���
8)�M�E3(׭�w���v;�l5��	͚�	��W�.t�F�$���F?��N��>�҆Q��f����nb�C���mp-�����e�O�duʆ��� 7�L l�u,F�^��ܱ��%�J�-U8�-"9� ����Q��bT��h�L�Gr
%�3�v��������gC�?J�=�X���J[��W�LH����cnޱ�/�8O&B�|��t�LRR�R�k�1T�|B�'�rmC�J&zz�d&r��#Ө<�}v>�i�@���+�]�p��D�W���Ŀ�Ui�N2��n^���]#!uåJV#�����b�����ޟ��w���G�a�m>\@��R��H���{מo�'>�_o������	���xϝ����Xn����5+���>�L�>��Ge;0'�6���3J�}�k�=���:�;�_qՉ����1�`�@*�ѕ�bnx©b�V�1�h�b���+��QM���E��*s����k��LJ)ժ����Fs]?Z�;��ÇS5p��M�!?x���hE��t�K"'su;;#Ԓ1�<�ٞcT
bn�u�bV�D�/��'�2[����2YК��"^��������B���U��o¨�6D��
�$-�Y,� ����c�8(ɳB:_��`#}�r�q6�p����;�J���P���}� �md�~֚W@���&�HSD�����bz  ���A�D>ŧ9�L��c�WZ��@�[\���UY��0v�I�a(�-YZ��a�{�0&��[��x�\D�p|�������1vb��*~��؆ ���:2�R�r��?
����v"7��\��7��]$�l>�˅��0b�>z�ǒ��W���J̫ ܶ����â��>�\�B"�(�$�"'f�; ��M
+J
D�]��-yM�i�Rc+��^O� �j�\�#@E�a�ItI�[w��>����}���$��_�,�ͅ�A��I���Ax�����C�ɭȮE�<a\��m=���Dm�F�簑�����(���f�y=�P��a�P.�М����fý��0x�D���)��X��pܮ�\iՌob ���w�9#�,��ܫ���JB��Й.��8t�R���dK?[��)g�C���Q�@nٜpWj|/A�XAjY����ϗ�����ݯT�kg�jtI4�f�L҆!�X�ʞh��y�y>I[ː#��m�%�c����R2 !uy��P���E�$��a��v,)��wH���{�g�gv�8��gC��8!�i�"F��1Q�}m�7d|y�F�l�j �����:h�@0@
?f�\K�~%�Y�V���ڊ�M���I]��)�t��:�i:�'��^�K�`1�f9����t�>h�H0^бcΗ��)��l��Cec��\G�2yԻ����ր��ƕ�c����G�N?�����E�x
jx�[�b©�8"�[�Ó=��-�Ŷo��z�����µ�>��L�6Y�aY�;�| p���'�}u��w��X�؜+��7.7��I������IJR�LW����k�G��'n��-D@�T	N����W�S�:�(�Ku�q!��
;���R(�7��(��1��ҬE#�]�i�3����Ibv�ob0|J^B,�F��u:�#w�����ֆ�ՠ�5�E�u�S6�7��sr��hˍ�z�A�A]�?L	)M	��pEN��J�k�'����X&]a϶��C��8���\�aF�s���w�)��B(�(a���D�β�=N2	��pk�}�zw8}9s��Vs�x�SM6���X�zwI��7����nr����H�7��/Nn��U�1�����I�su
��B犆�Pe�s�;�F>+�L�c�����A����,-'?/(�����y�eO�9�sgUi
�̾w�����[�Sx�3b���hw����	d�B݃W?ɭ�|��)�n-���lW���ԋ�cx5�Vwy�t`�g6���w��d���:C��G��8D�c� uA��B�1��
׬ޡ��<`�B��%:��5�
��L��C���rz;o��|���T��C��1��-�}�2�@����n�����.@����9�S~R.��,)F1P��Ջ��}V�Q�-��e!��E���150=Ѳp�%xoZKM����m����2]��a8)�{-jS��Џ�&V�/��4�?�R�)���ٗ�pKHP�<4�����1�|��VAQ�-��Ɲ�F�r��]5��{��{؁����2����[��Mj/�y��̧����JS���[l���r������%3E��i2W�뺒����s ,�l,`!�������Y�'na?��7!�s��,�7���G8jx�'����H�Ǧ�vg4�5�b�M|g�k��t��o"������<�N�Ue����%y[k���a�7�N�n���D��;����u��,+I9�Cv�s;fl�
7Q?��P��/�,�o׵E$�n&��Pڅח6(`�/;'ܞ�6�r�-f��*.q<CϟS쫍��j���%C��y����D��h������8�k������$�^'�خ�����3v ��Ī �Z �[�uv���D(��'�y���^���`� I�����*���/����u�����+t\���:�W�`�i�p�KET�Uv4\� f��ȹ����&� ���ԎL�UF]�������QW2�q�w~�``@�wK�9�'�m�PlάZ��P[�B���ܸ����ko�:��|��ZGqJpC
6kU�i�;[ܠL�)%��W8q�$r�H��O�.;���u�}�����]�gP�<|��ї㩫�:�M�3c����9y���N��v�-`?8�$U�e]i���q�y�_��[&�����p���`D���.��CP_+{�"︓�4/t�I1�a��d�T�(��3�������I�[h�㉠��+"M?�J{y-�M���ؒ��d�1pmN�z�#���(�E�=�yv������<Z������ވ��H��%��|"uQ�.���*��u��*���}.L��������u��_�j���L�WM��![>�\��T��?3�z����@%�(�s��K5�9���� ?*e�۴A��N��_�=ؓ;��"��"��������-�Z�l�$�K��b9��3�K_�>�G��
���Z�ʊi�6��t�̫��7�X?���D��όwNa�<�,��6�+>~�JIa�S{���֖U�J���#n!,!Ť��U����H���#._"�K��+�(�� �R���wo	�E[�z�/����5�B�
��-��IQ�H��|�	p*6ET�4���=����L���#�R�����S�7�vl��U��8K�����y_m�X�`����|U�9V��U�q��A��,F|`���] Xt1ٿ)�p6�o���iWC#���2i���%r�,��_D�g�v�ư��o�qI[�p�,�;t��r.k��/�()�Xz�v0���"�@s9\P��;����}X�^yIu�7W/䥘��n*��d��(%'��J���En���:#,܄�7{j;�*�vP�YnP&T���wM����+Tw��u��J�{�m��6sG���%ȣ��l+���A�jq���-�g��DBc7���,!�:�� �Պ��\{�r��SIO��
�O�lG3\$(�a2�p?o9���0����g�(�|LF� 8�׏���R�"`�=x��O��ɤ#���q �����힓�.k4����z�_�Ğ�<?*�*�gZ�:���hdl�8���;�d��I~a+��]���R���Tw��9 �T�v�X�z�������1��N��n�Y�Z���1V���F<�j)������;7�8�Y:�d�����%�~@q�͏ܯ[J䛷���M3{n�O����`�|h�W D�j �ǠoE !ꮻ�y�Zb�/�צZdUe�h/Gy��X�\�۲�`��~j��R�/�5ǀ7O)�U��u�z�r�(F��z�~��B�t�p��P^��Lui��/A�O�g��*`�?yN`I~�E���a���Ǻzj�0O�A����rX�j��~�ф
??��!?��D���W#�'Ek���wh�f�|W�p@��y�V-�%����Xw�[��l���`6�� < ��-%wUh�a�5�;b���
ǼPc�}M�V|��6��G�2f��H�X��Z��A0�Ũ����U� ,��%�\��å�����|_}.�VM�����Aֳ#�����27�j���%N��^��ظ�O%!�`���_�7��l�#�\���(�=upzZ�-n��z�B)VCF�Q���A�?�{;.���e�*Z������~���g:'")qԁ0�{��E6�$���g��LV����yѾ��U	�a���J��HU���p�0%���gǅ�W��o�{m�1�Y�X�V
C�ȍ�_kLp7�O��y��f��s��{ߕ5�2������f'E#JtK��-�zy����}/�k�#���x�lOI�A�3�U��O��s��/��߄����Y�6}h݋�U+dFŕC�6<��_��w���A���5���r�۪�:E$�*�TN��a��V�YSr�,
I:k�~`�\�m/�G�R�s��C@������?P��D���5�7�W[eO����
}V�͇�:�,h2:q�!�p�<�G?���#�@k��d�b>�V���o��#�)��K�i�g�+k�L,�YZ���p�����#>��L�,\D�K���+Te�sg��Վ�R*�"ڱ�L{ �K6�}�0#R��J�#,ȁi�a�2��YY�%e;�V~$HQ3L��������մ��?̮'U,��l6�{�}���-��k��9?p����⾙� ]�[��2m򩡋���Ϝע��.0!Ƭ6]�y�|��x|�;s{����@�ݳG�X}�lmm���/�?�VV��ȄT,��+5{\%7�2O��Y�HCs���1o�����e�m��������g܇�
�0�>!��+�����.�ֿN�A�l��V��-f9}�޲5�jy���*N98�&�մ�(���:��ݛ&�O�'U���O5���UK2�k�}�ckm�N汧���S�:����ax~5\c,���3��3vݍ���i�:3��jR�mA�Ô�_���܊��e
�+�ާ�+�>�6o��H
��������^+�TĐ��9���$�Y�<9�#��ռ�⎽q��{]Ⰹc����;���P`?ڽ��]�wpE�G�g�y�}~,+���&�Ť�7#x
:<����,�gDL�UP��7��? �GTV�H�[��֣7Ej#��"ǧ���=�(m��g��E��4�u�XZ��S$T��U��xE������� F���b�h������N�W
˙�9��_�P~U�qE��L�2��u@��;?ڶ���sL�@+��/�F�ʧ��9��?�bͬ}�`0���(������9P����d篇���4�mU��6�N��W��1�z&k�}T�$�|�Ţb�����"�	;0Yʷŷ��J\�3VЏ/)��Չ�=��@\rDk���E��ҏT��]d��7���7���yǶ�*��n����U��u���	�{CB�
�v��n
v�>D*�M^iH�o�`�"��n���{���=��ʖc8H"ɲ��N�I�����/��7��#{�T^�����h�ZL����%w��s���'��4�ƞxĩOj�Ԍ� LH_+I|n�u����jUÏ1�!��>�D��;��J��D�TU�aZ��5YtܕK���Z��f1�\M����>�@�~�3*N��ĸjk �p�蚋O���7��A%���`�k�Y�PWE�4��>�}jB,ݑf/g�Y]3{��v v�x15X�%wD�u�s�C��Э:h�|t04�\���p̓{<��N�A��lV 5a��z����^�9��
����Q$a��l���%���o!v�̝�Ĳb�7C�����(��R���	�'�f�;�Wy�N�:��,��k��mI\���{D4���'�������f�m�J2�P�u�yi݃��uB[Cϣ?�[b�? �H`ר ��(ɰ�D��>��e��r�
?�̓�>Ǘn�����]4b��2%Ѷ7a���q�ɫ���Z�SVwJ��^L� <J�*���_�VF��ID*.m�k��s6���m����_�+�6Г�
�+� �(�w˯��\)4����q�6��u���^J�td��V�)�'
�m:��â��m�����K��O��HW��ơշ� z"���a*�G��_p�Tj����>@�I����N�8�r���
�d{ӄ��7���o�f�4�PG[ܼ�w�w�h�N��׉��0
���v�b-�Hy�.1�2��VKt��8id��ÐU��2ƓW�3��՞�}���ݼgf��n[�(�U;x+n��7nr��:I8��@2}}��=�Es�Tm ��<���+!��s�*(�������|@���T���6:���4�����f�B˨ϛ�[�sk�����&�k�L�ƂP팟��"��)���ɼ:������#�l&�T3@��vޛ`��@��S��L��BI�+����V�_��9��r�L
3!�I��pr`�q�$����@�~�@���\��F��"c���Vؐ��N��!����0s�N� -�\��k��n)���Y����mIg�.�%yj�7o]P��S�O�s�W��o���6ӳ����L����5o�~�(�,H���"��F�?�)���	�@�^���`����
�LL��d�We��=-f����g�W�q��y��	f�
�	3[Z�K1C��b^ЃN��O�Jr�S͍����S����������71���Sņ���`P�\\�����[�$R���9���iA�g��Ȼ1U0fA�L�½�T8	S&�m�ƾ_��}o�p��H�����Ŝ�In�SS20�_gy3����\r����Y-� 	�+�{���yf�u������;�&F�5��]�]q��x�j���ࡦ��R0u##[H��}�y,~�8 �T>�w�[� �ᣘd��L��Y���N�hn��d�\��R2��H^�u���^ŵ����������{�y�����H�tpa���6L�FW��?�5��.�>��i�~r�
\/��M�����/�B������*��t]4��sh[�!��|���f�p��X���6�\�4>���ItnFѕ�h�o�c'<�9}��8�:�홞oB��]VG}��b��5����kՃ,Gnm���5GF
�D
 7�a�^����Uf�7s.�nz��T��,Y_K�Hm`���SCE���s�]l\5a8ReK��{�d�����1��4�H�4���#�@�}o52��<��������nL�i���O�"2v1�6ܱ@k���u����/c��y �\��Z�.ȟ~i_�wj�S��r3�?XH���Vn��GN��逿�MH�@�������cVͻ�j�}��,K�(��,t�h΂��<�� c��QіH}�hH��
(�l�Y��^Ry*X��jM�ⅡD��;�	/�6������� ���Y q��%O�2u\��������c��ql?�]i��4�u���h] W�g2_���[S��g��I�K#�_��O�lRKjeQ�=��0�f,��G`T��	���z2&T؛�1Tj	U�n'��1j`b7�� I��Gm�5u���B��>��LO�z.[u�ƾ���Hs�=�hġ�A�|��bY�̀�R�K�R��0���c���ŧ5�C��'� ?�����*���ꭅ��������2�ވ����[N�NN�X+{��솻�#0�����!�WT(��8�����Ĕ���i�vړ�Z���	b{���nf5Pe�qw�ip�X�)��v�ki�3����iT�V�P:@
T�b�Ou��P�n� M�q���x x��o߭��- ������frg�=��a"3��[���_�j��)\-%@�˭��}I�:i���qȘ��6�׶*3<��T}E@�xvzB��D4�삎o�*D~�;�f:�a-kZ�U#�Y���Vm�è-l�eޓ�\��>mԟ{�r�K֔��1��H5or|�ӫi��G��7;�����n1"��.�������Q�7'���K�xc�RhƝ�� �ۤ��)O��`-�
2�h�c�\�~[�S�D{��};�@�ϐ��շ��[C�M,��a�,&�}iA��d�!���_�)5��>�v`&;�,!ԥ ��e8H$�{�C^^7���G`ް�2�ec`˰RD(�r�T��vR�@	�F�w�fwkj��8�%
�p�� W<�F9�� i��`� jj)�r�H�}r��>X���Q��F7"3�a*=�Fh+��#*�w%�u1����?����%h�|�E��C�`/O����b�G�u��|��	KgEױN�qց�׌~5�^8���9�s"6�3g�>v�@�!6>"��l���R�\��s��&ϑ�g��*�)�CQ_W��D�X�AuW%�&�L%E�HlS����4����R�u���k%+X��֔X����xo+�Y�>;'C�Ȁ�J�˭p!G��B`;��p���Az����k��lt-�ޡ�viY�MǕ�=�����X��U*?�q2�ۿ����'uO�t��5�����wx��iloa�ѥ��L�P�'�BH��Kml%Kw�Jq0^�'
מ��Z�B˖��m��V�D������D�7+$.�ji�
c��Ų�X����ݙ*��ߜgB?J�9�B�:
 �?4���j{x'�E���K3�0�l��NU �Κ؎B}����.��Y��C�'��y'�3����n�0R��5U�e��y�,�������p�~/��576NM���a�����zp(��}��1�$�Yc}CUN�n����Қ�+/��m�B����3�e�L���}t����HQ����qjO�5�f� 	��W��-waWO�P������7����0����v��[�틀�{�S9�O�Z]��7{K��-|��	�3� KBYip $q�TS�@:��zL2� �V;f9w��;��o�7��4}��mjg*���k��TY�z݂}�_���)r��{w��J�!`T�f���tF�z�g�+��,>�N2��&("�l ^�ʍs�[��og�oЯO�����!�p��y(x">f�?	�[$�Z��눪�-T�GQ��u]U ������-v��W,������K������]#r S�7
!l�����'1 �a�����]�L{t�LS8�8��rL�2!ÒYO�x�`�؟W	��o�6ѓ*���0��-�;�Gp�M�����!C���wY�7 <����y��Bu���[�:ެ�b�����1r���i��1�#5.�|8��e=�W,��i�wt4Ѐu� ����A�4�s��'��_��e!��$��~RCRq\�@���MСS|�\%��mr�:E�i5�öA�A�c�X��!�p\���ŻT�iN5F�Ѩr��'$��Jv���z�����BaR���?̭�o4wV��ԇ�#�̚��"]#�JdAFx�?�ڂɖ���8ȳi
u�S����a+� [q�C�~�ѤC�ި������ia�?zx�!ȡX���ی?��
����W��t�_8�Rfp��?��V��|[��|t]돕���BS�CgX�5�[CW~�[N�GZ��w2�P��#�-��̓:(q�z�B�<���c��E4��{_�.ߐ��O�l��3aO�چf7�<U.z�<��K�H�:�GҴ��j��bȖ��WH�X���#Ԙ6���!,�0���Zr�i6Wz:��na�7�[��N����E�@j`���lV�*|_B|����V�t�V3�D����mKr�xQ)o����9i��Pbl�#��K��	��W�~�\x���ҹ�SI$" d�����SE�]j��X��$=Ȋs��e� 	�֟%�.�jd�Nʺ�������+ѐ�#�$�����@��<��`DQ��s�`�ek�5����g���Ò�r��4I�����p��E^b�Q�Kw�cv�PU�:v�i��%���e� ��w*W�si�W\�/�����X�w����{�utx�߁�P�rq��8o�l����M1�_��jCm{BZ|Z�Q�:,�A0���ôqf4��H7�:��kKW������P��8�e�;O�0�51~2�^5ж��	����\�pAc�q�'
�<<��p��V�����I�����M*���,lD)��6�F,�(K��/_��4�'^r�ѴN��vZ͔�� JMEDk�V�<L:����M$��'MN{ٙ]�/��H�4�9��&"}�|�?�Y=@�[�Wa��1Ӥ	w����FA��#� "̀)���(�ǈ��H��C(m��U����ǈ�o���Wvo�J������@�
�ag)6���i9܃4ho2l���8"�/'�5|��oJ���"�`��ti�s�+g�1�X��~�9�(`��'�����[}'z @�;���ݥBc��钙�M>��������]#�C��Wd݄�Hi��C� ����4�vA�M.��\�ِXf_�Ȝr��5�| �7�y�}�#�\��)[��R�t� ���f�e��e�<_2�e��zZђz��Pp�2�,�"���zĿk5{��2ͦ�� [g	��D*$�q� H��D���aU=Jqh�Drt �L@;L��E&8��E���-�#�59�)4�1�'��R�޹�����l��:�����ٶ���sY�9 �ؑ�3B�����]�?����A�������r��ͅm7�����. �\R�4c�l��󛜳���5UtzU{ a$V���]ć� ͂�q�q�T�ǫ���3o�To�Zd�n�v���z+�f������`#��	i5Ŏ�����ܳ�"$���*C1$W�5��w�Y��DV﫢Ü�=z���=�.��,�l�b�M��C69�S93�'u��J����5ؑ��t��P��Ta�a��Ih�����-��u��L��A3��~�e�j���7+���,z����ba���@R0�%{@��GP�.$�߸�Tv�
�g]��j�1�_s��"ݯϘ-�&�k�-�W�`"*=6C}�����Vx���������f���Ϙ�/ v����e�ߩ��8�!�ٵj���E�����0��|�++)����!d������E Ԕ��DU$��S~�����BN��k���u��?e0�rѨ���Dܩar����l7��y�==���%*R!]����v�#i�Ë��O�q��g��6�$8vA�[S��9qz����E���M� 50�/6t�I�|Bi�Ɔ�A>^�v7Ա��1���lu@]AG!q����3��qPK�݃I��M6��VX)��GB�e�C0sJf{����:��G�m-�͏�L�R�j����u�-X��V�&åPp\E+�(�F6X��iZ�  �A߀�3'6E��‭� ��cY����.+���塑�: t@I2����]�G\�?�
$хC����>'ح�"a��[�8�QA�i,��=��LZGʥ���C�&3����	��Sw*�h5#n�EJ��UM�~z�i�@(J[���Z+@5�|�
7J�S���ݜa�S[9�/c��Q��x��נ�~��hqMi4�Яu�.ʡR�c_��(V6��Ѩ��Л"�E#�������� ������;�ZJ�z��9l�Ht�0�h�UZ�iZ��v�m�x��T�bv����g^��`Ce��y��!�Ղ�rE��J�O�뽰��A	����)gϦ��� �)�C����/�}�%-�ɢ��^��(�kZS�Q�̢d[���L��B���3�aѯ:��c�.Q�{�+�w�>G���ҏ'E��rd�0P��)�mDf�����:�%�_�$6����YŒ�h��Mr5F�Y�3CN[��Q,��S�w�Á[�\D2��N� 4�Ԡ5��nwѐ=��s�i=���ס٫^�h�X]׏{���2�u�l�!4A��p�D\�	BP@ϮnP�!�Òq���_3�E26>զ���i��g2�ܬ�P�B�B�=�"����r)a &X[#�cR�Ȫ�k��H^Jۗ�T�%���@��~���s�%��K�ݭ���������ʛQ0�\"�I�8k��^Y�5�l���g+b�Ə4Bu�\P�.��5�֬�Kw2�?�8>}���2!l�G�y����v�iDB��sKʹЋ�
��A	�`H���hd�`��&�ܦY�Z��~D��L�z�3�~+��YJ�e��;՗t]��WKB\�LF�D���� �Mؘ2���Qgy��كr�M,ۺJEg~��dԠ�h��^�Y��nv��: ݭF�g���?/鹷���a�ee?=�Y�,�H� ?Eij�vP[��$ ���JI���E��n\��I1JyHªL�oҼZ� �z�+�MM�Rrp�����b�����#h�a�m��LF0�j�qO�F�5�����/�i_�S �4���������6�`�@=�)��������`@Mu9iFr1�YsW})�������M�.�a�k8s�{hߛ%� �;�}7����Ԥ��ģQ
�|�4��5�ZAo��(���'�tm��i����ܶ�Tt��M
*�-C)�]��CS���k)<xW|�:kdI�~伋�7,�&��{��̘5x2p�)hΕ`*�EX�����Qͮ��Գ sbU�9��9e5����7����}����v7f�v�)F��NWz�[�HW�v,r�6ϊ�R!�a�4�U�9�����ٮ�j���uU5�� ��B_M�%GQ[6MR��r>�o�C��0�8-�v��"�T�O|�~������#��ӝd�93d.��o�Y���ŗ���[:��5AY5��.�,�+؍~�lu3
P�h�K;f-��P%o0%����.l�MJ��	4������sIl�̚,OI@(����[lrJ�
����u����]'�5�^�t'mq~��|5���jB �����c�7�����a�����8�%��u�3U�tצX�E-���&I�Bci��īGr�����'	�W�V^�. zn�u���}����������ǹ�b���׳�eߍ_�u4[=2�%,�6sHs�o�\tN�}����e/'���y��#�hk,��%�9�,�G�T���S'���r�K�=�&�Ie�Nu���]�!B؇���L�hTH����&���������7f�ܯ4�d'��^]�5�v�=xhp�q��g�d��,�
_���S�;��(<q#���-��#x'�u�l;�A��r�4��nX��o1^ў��AWC����pxpMe� ��\{�+�(��k h��.���w�EB���AѡdSt�"��㉺��<Ρ�/M'�UUb�^�������!T����:�T�H۫�2;��"���1�?��F�8Um�1�!�^GZ�Dk^��I�3����?c@#�_�;�	G(o���8�9 `�r��$�M�pӷ=g��r��Qu��&݃�:@i�h��)�k}B��q��T� ��#JI�r�,R�ɬyA/��|3\����E�%����F�qy��������x�fT_0&e6���*6qA���I�p��8��\���D\_�u�����s>��jW�ˮD�1:vn��l�FV�,�p�4��$2vhjj���^�fۥ(�\%DE�����A{d2%s՟��y���M�_�q�dJGCG��%;�?��DC�M)c��mbx���xK�J����\���9���IOi-��6r*���}[�
0ef΂
�I�<��as���חS������|���2�6�7f��s��Ï�s�.�M�j'��O��И<U�Uc�j�t����U�q� �z�:�lK"�d ��k�]�3f;�?����uT��ޑ�j���:����t�*I9[�`��" eI�N)@1 U���9솗Ht������1�+�	!ԡz�W�ή�"��7ɓ-���q�RY���N�P�=lڛD��`����zx��ڀ��Tx�Jܜ�b�:>�Z����;ndݤ��ޡ<�Z�;�ǔ]6����W�݁Hco¢�W��W����Yy�@� E�@���y�G��f��`���3�ʆ�*��j�l���5� �>�*�5# ��<gJ��k�H��I���2����y�ц+��㫿�C��ړ�졒~F.xǁV��ơ.����+�5��B]���g�3(��ʜ0�4�p����}�2��P�A�㘝	���Hh��\�����t�%$v:J��In�|EjC&�6<j��/6t��Se�E�7�ěkаM��Ǫՠ�>�ϳ�-5w�kc�⍬�7P���seN~�΂c�.��44�'ee�<hD���b���B�^��z�/���~=�'w�	j���U�C�F�4�1;�\�癯� ��~]�$���)f�@%�B�[���ްC�Tl�=�E��k=�lD�ط�*� "oH��3*w]?Lgt��ګA�^���bX���]6�Z����5T�X�x��E����� YA����j����X�)�hl��B uV�8f�Q�VWj,���A|cmt�L��\=� �Q�������Ч󠓔���Ì߉�ܴ/Ǜ�5�J�l�"P#�I� �t�3sqO(���8J����l�M�d:�<�~M���� IG$�:>�������%!�ՒoYc������9�n2o�ڸ�4:�|1�tM:gU���$��w�J��u����?\�6R�e\i��ԥj���)�����yT�
i�ՃExj��atJj��������Y��PG�Ba"�"?�U$ԣh�Q��w��7��Cl٬�K�Np�-�;�UH�m+I������0�� ��I�-R�^};ɞG�	�/����_|@[K��ĸYe���qS��MS#򊗙0� ��-EO,w����Ri����t� ����{��Rљŏ�Mh�zI�r�=��ެU9{u$���mνe��pe��Xr=�y�ǡq��g��j�Q�U�Ϸ�H�,�j��zA�u;��\:�noeq���S��W���A�+)���"�Dya�a�j�v`;M�)�m����EZ��X��q���LRb�M�bB��dz[-z*3��*1gۖ`k��E�_1-�ie$h�Y�[X���J�1�G����ލj�xB5�b !�u��L����s����1&q�Aq�ҟs���Dtm�[�AI���"7 � Ȱ2>)�)۔��M%%�9�_�;j��C- ��)a�c�tԍgR�#n� �Se��A��U!=��8e��h�l���o��8��K�0!sgtIG���*1A���">|�ey��-��D3�* H쐯���M��@�_#�����Y�!�'�� x��ٛ�,U�����r
��<�dS��=f�@�C��B�/֓�[�P�~�р+8�ըR�8�C�[��x%�C�b`�x���6Y��p	8��k�����k�Up0/=��Q�W\������<h4�R������k�]���0)o�	�̉n�������V
���5$f�H�6T�������ݖWRȡ�:��Y�c�Og��
��~_\�Lj�"ށo>BG��18�(Y�;����A�w"�=����4r��2�XV1���>�x}RCn� ��h!ڵuh��s)�I��|�3e%�"T�>���I)���G���6��زq��v�D)�1�@E�tվ�3��`��ю�����1
�$��G�6�$�z�-�Ӯ���|��b^��d�0A���*}h:������E�f�'�i��=³���P^\ԥ�P�\�\U�P�*�-�b��#ަN����14ze����~��{�zZ&�(����M�D!�J@�%a^��L>Ɖ)s/�`
ڕ��U���[���$]|�Ni�t֔���sÁ�&��~:?< ��Uf����h-�>'j{<ٍ�lM�0�^ P����G��u:n�E٣�֏�E6�U��L��}ς�"���2�G4���v֐�T݀��ZGt�R5�[^��N��qj�M�f�k��s�������_���5>��d	 �5L�!��s��1�F �)�<�ȍ������d��M!��g��Q'^u�2I��%�%��	g����$$�O��2�ݾ������b�V6�XXU�T��N�l�Wr�8�*pƫ�F1���5a��S�x�+��KW��73��i��~%S���ϥ�bQ~+����c�� 7���n����^���S���UR~�T���Bka�#�i���1���'4�F��Q�T��P��ϔC��Y��8�]~a�]�`��Y1��V����M���0���Q�m���]H'1�	&}�����]���h�U�;b-�z�NI�H-yp��Hh��B�6��~c؀�����w*�o�`�8��v�_F�l�����?��� x����Тe��Mk��lZ��E�� ZBWBC�핈5�6��}��\�"�R}��\f���躥��V1�8+d-��tđ;Cu��5����BJ���nYJ�:C��F�>�J���Q��G�;dr^�Z��yB��?�,�&It���Q�����P:�keq6��Q���/�@��#��yop0y��+����,�S��hS&A��rXz���Dn�GY0"]��k3��#�0��o�k�qtٮE���䴲�#���LE��oO3����l��_�'������ٱ�J����j6�0�
 �AEJb�>b�u�y�w)�EVJ6z9�S�z�"�ֆ�8��������%[E��n�W�}g�%v���Gt��6����]AGzh,#���,8��{��]a�+lg����Gh�	�5(g��6�T�}2�N6E)��~����8$Ge���.� N��JR��9"=��Y�訆q�HQ��Yp�$[�hk;����&�J5�,ZpE�%%'�tx��?~0��6����]%h]����B@f�l�׎�JLp���i��I䈠��cTnO�XHr����7jE��b@df���n���х�7�C��>(���G>ښ'>�Dk8換��0����DT�8��f�_�j�<L/���m��v�˜��d��\�@�����o�R�� ��K�&�|��d�Ӟ��0��Bh\#=Esq3�uYZ6��ǰ�>��'g]6t~�ǅD�q1)G��U������:0��}��/&�/�"(�I<m� �H�;8�h����K3W�F�N��G����G�f�p�yq��(��JX����ph��KIh!���x�;�%��l�Ӓ춇W�`�0D��(	�4�q�h����R�|_��srE'����1�v@����⧉�߉1��y��'q�+����KEp����9����%�AY �Vy����&I�L9�H��lDퟫ*�ݽH����(x�+T6������>f��H��`�fL�U`�w�������4۸q�0��$*J~{��z�ǁ��W�S�/O�,��H
�݀��(�RK{�#� iv�w=�����x���O�t8=I�'���xI�������x�L\� �vH��^0�@���Z�t�⃜"�AK\KI����b!�*\���JL�)R���D停<8}z�]r/_`� ^ҫ�Ŏ�f�6���+�R�~as	�C��_����9W��8�*�pKzouW��)�w}U�^�{G}1	ᕪjFB�B�ה�&��RϕV�����g�K�Dk_��$W��9�@0w��L��<,�zƟ���0Ho++�91���.�dQ&�5X��f��T?S�<�B
��� �k�����G\9`\lݢ}C�rCO�J��U5�&�O�^}���g7
"��8�F�j��b�����*b��^I{1w��u
��O�5����6s�#܄{�7�;�-^~��iF���3����Z5Z������D�iz�'�΀��ԥѥ:�HmJ��b�c,��\��@9�g�e��bC�%��nϙ~?��*h���b[�$��~?���6�ݙ��{�IHb�Uy���T|�_���W߰*U���v��e��B��:f�.�gi���DQ���U���"G�ݩ�*�������±�@t�;{�� ꔙuv$��J9B��m���������60�%>���-�wFd� &�N2�j�&o^3���s�a���s ��jhT��LAy��.�Hx˝�F�Fj	˃�{�{UDӂR�^7���W���'{��o&%?uB��;����pk��U�X�����-�? �"��=��0셹h�-P���2Cf����Ն��a1�[�t�Ei����@v����$�"��m��������Y3�#5i��^��[� �7�kFG��e�/_�/�\� �v� K������%�|1`�����QP��bv��KE��."�W,HGTn�����@��B�IzR�"�4���R���Jm��s�Љ?���� �t������'�wyIcs!�9�p��ei��.<
��oU���/�?�Q�$ٮW�!����r}%��l����c!.�`.H�nj��qy{���zP�쉪���i���w����d�m��fxL�s�n{L_�����ϲMo	������U*@tx�^&�,�Y��d(¿hw��-�Aq���F�����3�_%r<'�fJ�P�� Ey�x���HK��TB�-c�X	�;}�(�d�\ ��NKP�d�R!���tOӂ;6e}` �#���;;�Ko�@6�Fz�\�ȐU�},�u�ص�83^�����k���GV�%�B����lV�䡂)�z��^=�V�
��,��)�':ŝ&�ڗq8��o�T=�0�o�0��$��P������{���d�Tg�J�?2�PR��+<��i��ə�=����ϛYJ��z ��ּq��	�4�{�]�RL�=k��Y��pv41����9��4Q�/�Ĕ�zQ��k��V���h?2J�Y o�z�T����cV8X��C�ZP���������kH�{�W�U�����ɮ�BzgO3�H6B�V��#�=T�����4	E�4� �{�;�I}�^�O�<�����6�H�5d���k Li����|M)�uV���Y���k%/���G��4���O|�sV���9�(�������Y��v�4�M'm�� �Bc.F{�Z��ʨ�A��/�E>�̭�XJw�w�{�O�J��,��Z3�m*�����������Jf 7k��/���}�߈�ӵ,\bEDe����3x,���<_��_�)�� �G�i�i6�v��s�@ϵ�esм��WJ맅&�v�@ӝ��V}y�����v�&����.�sP�� zJ~���/���F��#����tZ�٘��˶�h�
����y���Wn�J���P��x��"���QR�oA/İ�X8�D��wS+�u��O�?�����rN��}�P�;;�����m�|�@9ꣾ�3h�^Yd��u��.p'�0"IV��5?��M�Nq���#�xi�L���9Ռ�}9{g/��!� �����Q���#M�T5j�P�GU��4��׼$%�:�H��-5G�u�Ϛ*�_t������=a��pn��&1TU�&�cW%��_Uu�����o�qFY����~�4U3�5�V�iKDInL�jN�V�p���rt�7�˂�S��mA3�Դ��jZ*GJr�lZŬ�.�y�ƕ�"�O������Z��Vo�Q9�o����~�� �bF����T�ͼ�f�PtL�:�;�L�ڍ��c���(LQeY} �uu9sΡ��[��;�6�b��$��]��әq'c<1��靅>�}~x��i7j��;'7Ѷ�����#�㕦�,�I�C_�ۡ��!0@�m|H��\#���εj�� "��ߞ��y��F�/�e	}�*�s��j��s��,a��m�^D�P�r�t<
_<��2h��M3�7 ��hb]ў�a՗`�����ײ����"��4&��IeE�V��C�5,{8B�FɂAFN�~�/O�d��C�rաK��n�̫�U���#z+���|p[��d�d�A"`���e]Hn ��й E��֢K��	�z�cqh|Wq|�������iDP�M)�Ð�f ɱT�!>c���3ڬcS� �v���$�.�����.ԧ�m� ,Q0�#���,[��V���lL� ����߭�O���&.c�ꮨm������+
���B�	J�����%��d�P����l��W�$����2�m]�F��fͫQ�e�Z���ܚ�D��QW$naY\f����Yyog�g"�(�����b�!�D�����60ƅB�n���>�@*��G\n+�(�BԮ3����ʠ_��zX�/:���\�H3�{֌�×��Sr��uq�����5#�<��Q����Q�G|��{��:wu�͛����>�� �d��Q��)z@ʄd�Bi�G��r�=�����h���rFc�F��F�.������ aN�cP�2�	���;x�<��(�q���1a�G��\�B٣���+f�_�4�ҾL?��X~��^mR�y�x�
nIH�4�z�>�YTإ��Q ����_�H~��٘Ӂ+�>���^�,�oo�#�e�i��ߓ�n�h���G��B���8�>��bA@*օk?�(�N[�ʢK~��H0�ˑ��UL{���q��)�������K���d�ôa8�}+S��m �$����hsE.$g�g��e��-U[/��&��A����a�R�2EU�jl�G�^�.H�A9���Jd��s�ڳ��
k)8�x��b���f\(b��w�'!Ou�Dy�S�T�?L;�q���V�X���#��J�5��1HDJ6?�8Y⏜�]A(�W%,��⎸]��b�_.]���@P�aR���w��Fc����C_j�*8�D�L��AdTzf>���,γ{�F�C>�R�J<�mr`�?��X���Lt��Q�� ���]�w����N�ɥ�>\�٩�'�O+��z��ߔ���]��c}G�J��E� KC��/���^苶`���t����!&�7o`��M~h�~J��8�&R�����Z#���w./���g�H�^#=��Hv���-��<���Z���HްL��<i<�Z
�
��$C�X)�;���U�~ދ=ַ;�he��nl���/
%`�c��27d!���Y��b�K�'�s��w��45��/&F�3`�&s���5@��M�`�S�K��ƦLN����0Z7������� �~�DJ��)2�V*�&[(��zY�W�<�H��2��`��:$�Em(��6cO����s`�F��z���A�/>��%�[&!�A>t!�9M���.5�E��сA�w�B:��oY�	΁�'f1����nz�	~����%�D�?ZEF���-��m��X.��b<��<(C���&k��s����jb�ҠY�I~�_j�L�Fe4,vV"�쩶��@H�G��Y��������M�`O�'ɼ�;�f���~*5�,%�LX��m7K��E�ר5��o�iG���9A�D�����[���آ,09�-���8Y���'%@�B;��Ӭ5f
�#)��ٜu[��)h3��B�a"h��02�U%�x�p:��n^[-y㚗cD=Ǝ�4��X��-�M���:��R���1hDW+OUBT�{vnC����6(1\7_���B� j�b��ϫ
G�ٴ0ET�U�U)e���Y1O�G���p��X�e�bz�NsV�S���[>��?���0V�.�OHQ��D1 RI<��}��f�8v��3w�M�{&o�6�aA��lt��q�?Zl�j#>�b�C�*��u*�p�e�f�do��c���W���m��"��gֹ��� ������q�,J��c���ٯ]9Q��QK-�T�_NO�;����➋�8=�i�ʛo��.> k��'Pkә�g܈�6	rk�s�$�b��ETi����d�:&xej�����9�(�~HWx�����<���L�W9*�0�[��7��������4m6�Ѧ9�B����������-�D��n�̟E����-��T���M�F��q[�B�_�)�A�c"r���N�6���<5N���ɘ�&SI��OfW�x��Q�����3x��(�5qb�O�c���Vy	�IbcTo�����C7?�P*$ X�QP�28��h8�����v�>��(G�ԥ~�3O_����-�_�J氖z�����װ9RA�)�§V��s�1�#4ǒ���FR@>��M F�a+�F�J7k��s3�hϥ{Ϣ�f�����Ȳs)ص'Y;/�0M�Y�Ý��u� ߸�2ǥJކ��/Ę56�ꡚ�|���M6���~���A�Q�e�È¤� s��2�3^J�3>�h�[�����-
�q��=���GXaPÜ������%-��.ʬ"��V���F�N��]P���mM�8�8��mǲC��Bd���<7��"��E�ک�IjO���jf�Ά������{�r}��=9�.IOKt>���r&���t���p�>�Һ�m^Y!Я�GdS��]�eZ��Z��>W�-_}�bM[��s������� Z�. %@�{�9������x+*� +:�g�!B�Up!J�Mڍ:ЩJy3�:e:��aQ����ıK��j�'�cb
����_m�)�T��/��wU��V��=};������S��K��d�
�?]����P����2�N�����C���gR���A{��J�w�L˷1�7�+!h�"SF/vsK�=���U%�c�W��-/>t��Rwi@i�z���ud��ǡo$I�}�	���P��屵�J�qAP=�	��c1�1��ې��_%�����u��k����![���b����N,I�O:�Ku���IW\Wa:���'"���O���u|,f�����f��ݖ)�]Z(I��q��0�G��n*1��tk��L0�z�5Y�@�6=���釘m�5a ������s�Z�ϥ��q��w�̩!2��m�|AInq����:�����W�^�c1 ��Ύ;\�S/�^_��A4=u��S`�(��%$d8���/){��~���w�߀��5��o\���đF������C�rԿ��@�sޱ�w��qr/��k��N�'ֿ�O�њ�X�k�̙��m�'��S�
<T�şh�c�zp��[4,���q�T�����M�A�J�x]}��g4� ����0e�H��N� (�~�|��ZGA��fZ�|�Ԙ�0	����3$���������5�A���.,�rD�9Y��%Y�V�(�I(�[[��O:��|F+!)o�Wu�ᖟ�t���;�`V�Û;�$$��_�oua�n��2��A��'�Qv�C�C�O�R�.͝Ox߫��!�w����>��lg�n��.����N~W�F.��?'_g�63=z��	~������0C�fK����ˍ����ţ�=����h{��RFVAa��P����g���Ίg��1�b�%���5�9��d �u��)�k�⼨��$��2n�a$"<a6Э
��dT�d�ݕKQ��g<���Q�]W��I ����Z{���y�C�}����NS�V譵t�<%5�\%>�I��	C����>����ǖ��R��Zv��M&F��E$�A��Ed��`����y������}���O�s	.^� ��3_C�9��:�7���W�i�쇥%�+F7�nֶ��H�I�!r\���b73S��9�S�_��biM���s�C�hZH��u�#1X�K��~�YA��M6?�U����G.�<�����f���q.�T��Y�[�V���9����K��5���1��xר���E_��102	o�ԙB��������Mj�<�R8<�3�S�i�q����H|A�	�����o��2K7�� sU#%�}���Ds������7f}��B�#��0�(Q@(ێ���P��Ɠ%g�y.�G���H�fԗ0	�ɮ3��&�3�f%4�U�7����o ��쓥�ߞ<���Y5��[�r�If`|�Y���e��b�3�D�b�mmtdDɇ}��!������"��5��K(8����)-y#��-��hzv�Qtm�|���]����*�HP����?͛1����M���[��C�֤�:R1T�Xu�xp�װ�g�ʁ�(�*9�y���y&	����$y��I���rϘ0sD�6(��$:l�z6B���ބh�1�b��5��W��-�.H�w�]cĄ� �/O:j��?���a�Í�^���O~ڡ�s%�[�[=��|��^�������QY8od�=�c��b���v＊�U�L�8sh���5_h�V(�����CP(�В
z/�}�8��v��(�=���0�Fj��-���x"=�������0�)��]S�d"˵����I+Y�����ɇ������1/�������_c�.h0N;3�l�/��0s�e����+4 ��4ŕ!�h� 	�����g"h��^���JT�S�(Vt���$��V&][�"���60~��j@[�ͦ��'�թV���[I��d��m��	�e�j�k���*�� �F��q�����\��@T$�����\}~���"�'�V�P�Ht����+�`�!���Q���b�Z��r>�1�A�版�Qgw�	�?!S��������^�nI$ǹ�X��XǧQ����@I����-U8�Zl�\&��G�K��=��$:Kz@��&R��<�42)-z�������_Qfi�Ђ,�������A��b<䪈�d���;�LJ�*�0C�e+��D�q#�b��������~�l��4zb����e�l�����n����k�DC|%��*�ib����+�6j��`*hAF�Mp:������ŝ���G�L���+s��3�=��o�#�L���A]�� `7��ŝG!��m�������MD�Ԫpx�h�pɭU�9]o^�:ĖBBW���&+���k�>�Ȍ,�Z��U�<�X,���
l�f�AA�ǃ�A���nϕ�3��Dz�4qr� �2R�v5��v�qd��u����TCj;���#�$yVׁ_)�ܟUK�ZQO�x\�ި05�����k6��tYmQ�P�l���KʗI,�(��C�<c�R��g&G"EӰ�a$"�	�3b �Q:Ϙ�*�]E�\�#�M�BCЪ�y3$f�tn'��^W����e����`�j�K�ʶ4=�L�a5��Ւ;\��:o��2vW��{R�
�X_?cj�}��Ml,Z��׾^R����!�I']£��J
~�8	BH%C!Ue�~�llD0>NV�ɩ��芽#�BӁ`�||�[V��0@jSQ%�b�c@߷�}�!������!��U��G�^�4}�]�?����왩R[d9�8�x��lЅ�)A]��s�[�(�,�Cr�JIq�2�?m�pQOT_cG�ps,���=>>����W0f�6eM�~sKB�ޣ[oW̒�(�clX���������d=��o�2D�ͯ|"Q��V���q��`�YKw�PP�Ҧ��阧��	�TE�A�(F*��~���.t)>��CS�����m*O�����~�P���p�P<�#�T�����LD��b5dm��c�\������Q���myw�=��w�<�����ko�#��Bv��QY&�_�G�d\$�NvD��:�)�a�ʤ�[*o� 7϶Q��۔��.�&FjϷ�������Jv��.z!�p�-�<������X����n�>��
8$�bQ�1����R�|T`9�7{�sE����	���Y3��Z:�L&L��ApUB01ˢ�k��	<�f�pK<�!���;E��ܵ�76OϊO��=re�}�I�������I9΄n��NZ���r����&���i�^4�Y|�i��K2�Kk�B/��8 ���7CQAK�A����U7�k��e�9�G���;��+��8���Dz{�P_Wd疍��LW����0�u�q�K����f��4Y���1��!�;�	�� Yrw'�3X:-�c*0V���� H��<1�{Z���_�pQ3�+;��?o ��>��( ����#f-�ܳl���e�{qFp�c����U�PF~r��Sk�ȐK��A�{��q�'-}2C��w#zC�6��$��0��$67-��Sh%�9��?��m���KD�8+�m�X�9�|i�FOIO��O(l�!|����Q�`}<���'��0��v�\;+��T�������s��O���u>ʠ��T�R!/���H\Q��+ɋ
Kn�{sxxo�rR>[v;�t�K�N���-Tǔ�����iXa_�8v_���/�)���hm2t�7F9�b�p�o��^qG�]Dy�jF^K7�K`SH�SP��xl)
T�}�8S'�_���`N_z�%�U /��ug;N�ƿ������c�ꒇpI����>��� f��y
@{X�$.7V$�ҴI@E��M!�[���^b�h��T�� �-	haB�Q�QB�H�z�LP��ȃ�D�q�.]U�&��2��#Ёٍt@�f�aT'Y"��hU�12�:���j�SC9a��in��l.}�Z�8ݳ�x�n1�WÏ��b��jh���dy�m��N[L�Bp���G�0曃aK:;#�/�aّ�F!R�����(5L/���$Kq���A$�:���/YB���6y�:����0(y����P�����WpG���D��~��r��C�����r�ף����!�� ��!bg����F��z��. �\s�E�B�4��@P�O��B8`�n�5�&�Xߛ)�Dw6��:�m�x�*pzO�|L'b�P��d&AR�"}��v=(���qe�o!ܚS3�Q��EEx�� (��aug�xeEɼ|ی5w��A�J���C�ɲ┼�(��S�h������I�|hc���j6n�������B���>�{󠌏��^;�q��V]��ތ���"�]���tR��7�:�E��p%ų�s��!��-�_����+O�1�;[���'B���F��X�Ui)�._�`Ј=!����n�A�L88��&�'%FHEI����9�y�M%5�4�n�#���o�"R2N�&{rҡpYPVR��T�de����ڭ�tĵ���'XŠ�:����tn��ie�3�[
���?'8��DP���_*��h�N19��T�TPR��̀J�����ЙI��p��	J�uce=���QP�j�-�+e����S����q��aYw�u�T��lt�R�q7d�H��s�Z�Pvϼ� b'��^o*�pÌGZ�\P�wy���x*���s��/ytQknّ^�4�s�_f6���Y.Ħ��@
x�C�b��={&�o,=��]��+�2��/�;>�Lg�
�((�=�Ӹ�� ^K�2���L��#���m�oϒ�zxV��j���&�s�NS�����2@c��)��v��/�w�	}��,�ӵv���2i�s�޻wU�"�I��^V��ۡ3��
�h��?SIá\�߿te�
�̺�_�795jR\N��_*�%�-�Ӥd�(U�1�V<T����c%!d?�)�W8wF��=.3����.�`p���o-��w������@�ӈi);~���|d���n�(��"��1	b�1�{�@Gֺ��1��]��86o��$��Ǒ"� ��X��@��:b�,_��Z�[�4�	��5�� ��kJzIfDνG��`��	wkrkù��ד� �3�|������Σ����c�8�n��o��9�b;���&���k�+�c��҈�O#F��.��~u�_����OR/1m��H��wՍ��Q����`稚�9��E���;�շ/�ƪ��U����#������
��7�$0V�/}�"P����E!�O��n@�pg-���6����Ou�;M�Vm��T�iJS%3�Cf��ũW{ڐ�,~ų�����}1%��z�3�Nxݙ�h��9�)�|�t|�eً	�nu�ng��2�H�s֕��Ȳ��Ԟ懈�2Ph�nj���#=A��Z�n�!�M�����Q;���C+�1�LܑkKB<�)��=l_�`���Br�n��YS�|����[$/�<
V��8x��#j8v�6�Bl=b�6nU�P\^�
zB��U,�i=���Y+�s.sbЅm��m���L멄j��$��Oh��$�*&��E0}Y^f���N�+?�����F%�uH��N���p���g��ӕ.��Jn=��e�7���*UI}L@r)�tu9��?��D�-�&���3��{�˶��9����p�(aâ�����{��_N �%lI���D�}���`~4�F/�Y�WJ?�3D�����b����.�vK���8�N3�泩&��}y���l��F��'n�Κ����F�͊uߴ��"Z??�c��X��
��j0�/B+���,����sm!	&�V�Wv�De'��[W�EʪNP�`h:N�����o��,�MU��)4���`��+�����f�@��M���!? f��D���r����������R]W�x��;���|�������-DK�������8'	�@���
��0�h=
WiT��,��"A����1��H�\ǝ
С�/S�x�Z��cW�h�s��W�08o{[P#���L?�7���t�>Ʈ0��������w��!Q
Tz���y����0d�Y,Y�<��~/J�y$��B�t%�#*㽯6�fz��Ҍ֡����j�q�j#8z1�Y��1���OXz�>�@�+�4����Ŕ$���m�BvMB��`���rL�T9�|43���T��s�W�̦�!�W^)Oߐ�Ǽ+*i�Qק�������A��{��[��Xz�[E�N�:
��4A�yy�]���Pۛ&�z!�
���|8��LmnF��#�U��/")�8{g����i	:|�I��{VZْ.
�AC�Ӟ�SFQM/�.��ˏo�8ɼ���!���4Z��xl����Q�57sG� >{�}1�LK6A�='8A�T3:�ڧOVbZ�5�X"L�:l�"���N�~A��!� �?��:���
#zIM5ZiH�t�4��K�ƶk�i�i��Ŭ���|y��Iw�����?�F$xˈ�O97��&z��M/.��
a�p;�(���I�OG��1��o!����sؚur�S5c��k�f]�+�z��8V	u
q�Q��9�j�p�[~�������|?��>�r���4���ͤn;���X�����<4�
U��(s�ċk��X�S�rK�eEUaA���P+�)��BЇ����z��1q��2r��̴ƈng��>q"��y����Z�(HI�+�x�=	��ߞ��ݳi�"}�G}f��G��qh!Y�������E? ����y�0�;���ҩ�Hb�n7��
ܛ}WmEU�ᒟ���F�����s�Zu��k�~��F��IvZ��% �������H�=�t%{����B˨�Y�"�e��!�*0���B�+�����*��� [
� D��x x�wIG_�����iS̽�7�i�OG}���Y�qL|,���T����iQ��CH��:gN�U?Pë"խ۩�s�Д;w@3��{�DrbN�8���/7�� ��s��`K��D��pI��[����[�o���=��vK��r��cˆ���&�v7s�����,�LH��i�+H������Q|%�,D����g�N,QYe�b����}�$T�Ti2�|���@���j暀��~k���+��7���Ew��z8O�T@�<�3JiWh\Iq���I�c���r�Ʀx�!��lF���q�ޔ`)>,��w�PV�T�o�p#����jE�������gb~�4���P �W�8�-��J�y�Д�Xa���rrc�<
���
�[��Q��44��7�w��:�W�@1�t\���$�f(���L���i7�.E9d��-I�����1Ɏ#K�)�:����8�[�7K %�i��tuR��Du��%��PF�0v�,�@��Y��r�=VZL�����ſ!$Ӓ�_��f���A�ޠ
����^NH�u!��E2{���$H��+��ʉ�: X[���.����i�ƦDY>рD}9ƴ�E�L%� �5G��H� eݜ��L��v{N�Ԩ:Ul������-�4�P�N�&]#M�OZ��/�dB��6d�����i�
oOE�j�=/�P��&f��~xh���W#>��Bn�TO
�~C_D.r:I#^\~&���h��56Z�TK�ު���ߟ �`��19�h��<b.h��������&8L4i��"�*���g���	��ӂB�)0f4{����٤T�	�xk�h�ј��:��U��T�{t���ϛhd"k�T\��ןQ0�aO�����H<���>oߗE8�Wfx+�����#�B�(V�P�H�߱R�̸��Be�)�\H�F[��"�P��W��7֏��
m~��b��M��F�E�
�ŉ$��V���������,`�a�`��ϳC���Ǜ����:|�*,+�a|Ԍ��jDTl���X~+s��1�4���
7t�~�4�?MZ�ID�`|�撹�]�j��'�.C�T���O
y�N:õ����ڕ����p�'��\���Ad��@����W����]�@�l6����ż)��q��HYe:�'���?��W��V���-e/�}����4��e�|��_�}2�l���u���Ho^����
O͛���?vƅR�S�n���k�C
GO�k'c@�4�}A05թ:=tߌvp�;6��l�zk���}XTiM����F�1���eb�e���I�v˽1u�H��w(�(��{�{t�`�,5�B�7�2D;�"�ٌ��>?�� �sa�S���1���h�9�"�Z�n�[��g6�g��G�蔺��� 1M⳹�Y~��v�Cm�Y4���{`J)bم�.r�&g�)�l��;�N�f�*�Z�ɥ�O��j�?CNO��^;�(���w���rtG��ܽ�!	��]��g�����O'���o�v�{��q[� -M��K����ve'U��$<H3���k~��?'��M M�O�?�]n'�* �ڷS��2�mBza(C1u�v0^�)�Hz͘��:�b��X�<�������*`V�l;PL�L��ї�ʂ���6�K�Qc�~�� ~ŠeD/�.�AP�7��Q�՚et�=�|L�ʕ��I=��I�t�Qk��_�B�"�(�,e��*D�V��Y���ٴ��r�eF:ދ��ga�V�L�MZ%����ج�$����[�����}�CZW\d����r��ĥy�'�-�v��b��eF;>�V����TV��J������lt4ՙ���O~>k�/r��I��{�n���.4xK��Vi�hymQz<�Jz���D3��?%W,Z:�ڳ%�ew#*N�j�~���o��/�gҼ#��5���v�*����oz\&�pn��	��*�"��r3F_��z��
y����I����熄�e��oB�/�0(P����'�/ �$Jc�Z��j='���F������������*�0�&�3y��W�g��"���m�T��fN����*%�VW�W���oa�9"�A��a��C�e����`�.�q{��y��g���z��M�^�$O�V��݋�����8�b0�;�Vr��u��UPj�!����=JY�2�H!M����#���F��tR�`����7�;g�v3]��_r�j��`n��9��}�Y����&�J��iFʕ�"���,\�T������q5�a�i!�Ԝ�s�pl!�m{�F��F�:��&M|�Lj����i�Ƀtsw[���LyFEꁠ�i�E�$�"h�0�� ��S��V��aɷ��%��B�>賆������8wO9�ˢ��T�����uZ�<m�>�MqgW&�$`mP���:�\��"1"��4$7���y�	z���W���롯�IQ`�R��Mń� p�`\TSQ8����ށ2@�n 0^L֔G�~g��︶�������hN`5�)?�n�ktJ���vǐ�X_�?�wj�ϲ�M���yz���6����%����BjVǼ(�0�#ϙO�Dx¡шD�� �VT�����`i�Œ�0��ay96����,��Ge�R2f!ȷit��b'�p>�/��r��3��h�����k-=e�����[��58�T��.O��!{X'P�o�a�q�4�����{�p�%k�N,�_��\�ޫE?X�@~�y@v��E�?���`|�����{��뇍��n�p�Ej�}�������!%="��Z�A�4��S�r^n��F�~�qY[�?ʄ��ΎS@嗩7m�D���@
�w:����H����{&n:KH�d[�������ݣ��S��e&��h-?�U	����՛`����d�>_M�VY�:d��g�3B �kCXj����(����F���� �� ��_<��/�o�=f.
�26n���B��v���p��4���N�.���N7���d�����+d�sUI�ݰ���CD;�\�|*����oͷ�^���r����jhiI��ms[��pAD��~V���� �JdbSg�v���Z8u���tN�o�K�|�S�2bl[G�#�����W��yq��"��0!�o2���&	2�M��sF,h��9ݳ9�s*����ݶ��Aν�I��p�����W�(��:��|?�q1����I�e�74�9�\�U�#����8r��H��˦�W���x�U�;��U������� ���|+�i%�!L�s�)X�!{ϣ�¬7�S@�~E��Bk�?���o���,���p��{��R�U�q�Jb��	@���#�aw�S�����:	ebP��� �{N��nx�n:�����;m]~��A�^7;�
֩Nv��'mfʺ	���)�(a0�+��%%B�8ŹϢn��Ԫɉ�29;�	���?�~d�eT=�2����خ�K�3OӚ��Ƙ�@i�2v8���ai��GSY�vw��)�=;^���!�,M�܀Í���%!j�B�q�����m9�8��iq=n��)?��ĶL3��9�XB8�-�g3�E�z�	�T�^R:��؁�����2��I��M�
3~��Rd�>����HU+������E�1�����d�'��7%�z�mh�7 ���
�8�`�w��Դv���I�5�)e�^��mK��%���4��hl��ȷ�3�z�~����m��¼�����"��A���O*ˤ�yWh
��������I��,BM�6�{!7
o��e�����工f+K{�d�:��jhU;n�K������3�I�EZ7z��oMV�GD{U�=Pʸ�z� ����j�}�<�%(���;Ր�c����\`�a�̟�, R8���B�H�S����æ#\�n������:_��(�Z"�U�q�����q���҂�6�V'��;g�#�s�x�k�/p��FcE�^.����B.W�-���|�^�$N�.�vl$�⿫�n� =�x.f`0�Ex�
>�pK�9"�g##�Z=R�y�[.�=��6I	"��,�32lߝ�jj�ړ	V�եW~<�w��[FoeaЛlZW�b�yn��:!�Ea�1&������}܌�y�j	�w�+�px;-|%�;T"ݨ��E��uc�]Ͷ � 1��>�5�m�z�ȅ2�
>ޒ����
	hC���×�?UXw#c�
9���m��W飽��3�	,	W���NPɄ��#U�o�G�� ���	&DZ�$[W�^�����P-7�N��ٗ� ?�9��?�Y,5���}r�������-ѫ:�G>F\W��j�@��Z��#r��#��la��G��ɋGމ��$��keK8!��X��q:����bE��9,`.&I)?Ҫˑ�sݏhK�5\M�g�|�E�U$9'4�6�S��m\��	�L>`
^jT�}�V#���1�2F����J%�;��~+�3sJ�
�f7�j6yJ��=ZI/[�����*Pg]U��
O�:'��JRA��E�Q�,T���S5!����y�A�"y�����(z3vY�i�0T���6p_:��3Z@W�@y��qp\!F�j�
��P2_Tx́!�� �埽G�K�llGjU��e{×��8�Oi_�\�|��M��J��B�h����G	����=]%�	��֯��{L�`��:K�>J�8i_עWS���w�V�b��k?$�7����G�0��@Ձll��@�����5t�~;�5�Z��#����1����9��$M2�\���jY����;�	7A��	�BLF޸���;�1�\���ù3�mٌ�rP����ʦW�9G��{a8��o�Y����8�t�^��,�_
��_ί"ݦ,��(��?����4ϻ����
'�GRIđ<�\#��h <+�3���1+H�(��"� s���T>��?�0_�EҫE�L�D	�M�"�����bIl�
������J�
㎎�-��#�3����7������&B�3dCK��p��tm��Lя#֐��|�����{�1�yظ=WJo�������U�!oV�$йy�>)��w���]m���g�����,P�t�����͎L��y��Y!@���I��A��26d�8Ki�T3�/�`��a��&U?h���آb��󋁈x���(��@�B�y��y�ҋ�f:l�C���T�'^-�m�j:G��ӧ�@LԞJ�ʭ����d�c��b��p]��y����ĝ�@(��;r!}�e$0��-��K�ߔ�{���#I%d�9����Sq�t�vz�A:8��w���UZEg���A^~|J褶tr�9�oi�`,��,�$���x�^c��{x���`Yd����H���g
{r E�����X��$7�J��k�q� �hc��:+�N�h�����Y@_�6L4���K|�yP�T�>l�%ZL��e��9�L��$��BJ;�%��v���a��������Z[�v�-׊#)ۿ�4��_N�Y�Rj3&�a���S3�c3 t �;���鵕a�RX$�h��n�����~�`6��=��k�Z�����슊Ő2� >z�� �?2��UvG�%T�����ܿ���?��S��f�׹�bgU?}�6�ٌok>aF�wW7`�Ie_(AE�Z�)�@،/?g#�.-	�#�T����Wx]m��C�q�.�(Ty>,���p�MM�6���V\y��hx�Ϗ��Uga�?"EB���QE��� 3��;PcO�\�6\�����c?�x�h?㸊%��z�]jX`Ɣc����q�>�$��ŋ
�F�NƖ�.�PV��
.�2ʑ@�����.�6S�6'�����=����(�SIﷇ��<����B$Of��4�6p�a᰾�DFc�]Jx���$���V�6���Sb�KJ��&fig�%�wk�n�ob���Y��e�+��ޚ�����2ƯF����,=F�7�,g̓/v�@b�!|�}��N�Ha����2.t�k�����9zEa��Y�PQf���6.Gn�q�x#��4��J���;��ݫ~?WX��5o
����Zz��y����f�̿�s��X��Q�^;�`1����_Lb��X�ϸ	��ځ2�%�����b�eU�]7��g *�A�����At�L�P
��;d�C��"��,�FT��%����x?.���j'�,�0wQ����������U����j*�Q,W}�?�L�������s@�W���(�X���|�:��ù��H�ǋF�����k���)˸�cػ?��D�]��K��)���_������Ʃk�\
�4�ě�<�77U
��� �"�c�,�^���� ����J��+˶�ut'��f���Ֆ�����U��_��8��^8�6�B���<��.�h2�.�*4(O�+�R�ܬ�G�y����G�����e!<�٧��I��L/g�䔍��H<╌�?'�d�* �H+fё�b.y�wn��<@��!7L]�������3�Mw��k��0_�詔^��ɢ4�q~R@��ul��(Q�i�^���wRǏ7�?
�%��+ڎ��h7��&}��SЍ&��z��&T������6ai�?��Sd���6H����{��C��� �yGm5d����}:Lv1�3�Kk�e��_����Mw���q2�E�J
I�&7jr��5��<�8�b��nVI=}`����~`61�J�0���^����5Wk.8��<�io>���Yq�0S"���X�e{o��:���ߣ�o��>� \�J�����z�����T��[W�d��O��Tt.�亻�@�#3.1��v�L|���pr���"5H�5S�}-��|�۸�2��?{�%�V)=6��׏�2���.H�o3���?�h�E�*x`�������[��zG>�3����Of�rw~�bFS�q#��=2��.f��;WK�ZW�0�&Q>�x{��F�V��ޚ�j�j�f���U
������1tjÛ%��ˌ����v�|%��R"���	%�c��Ƃ��ȭ���0��B8�b�}�CdR!�V@Ăl��)�A;�=
�d����1�Y�5����y?[^S�.CXӑ;h�I��`��Z���m��v7`�=�t�^)���m��v�����.W-b��\LmA��#"U�F��� �@�CV
�p{��O�f�=yߩ�4객���L�-�����	yȢ�m
j_��P\+b���'� �8�H���Sm����&�\��uB�'���� ���4�j"�=6�'I^��-}�j�|՗�
�m����(�ݶ*m���}��/� t9�W�K�L-���,���Ѕ��]��#|Ԡ���K�
^��δ>N�p���&������.F�u�:����w�;�gAcf���S
��&ŝ�
̣��|�f�ȼrcQ���У�ڧ( �V��S�E��C�x�V�h�}�hu�,yYN߻!$�i�:/s棳��G�0�ʰdp'�em3��-�di�e,��(���z+Ĺ�K�N�e0���с����=j��m�J��Vܽ1D���?V��_����1 ��g�B���PE(X���?ɤ/Ӫh�"�)	��Tk�2���C����*6�Ǹ��J/'�+�j���Lf��XIk�
������*<���ӨDN�H	��t���%>ti*T8�8P񢳻g`K��nK���s��a�n����)�O�N	�ѻ�}ي�F7����'��p�'Q��s���V�.�n��;cX~^�����-qƾB�l���|?xI��c�IH]Π�9NxR�@m\{3�ό����C�;ȡ8_���_
�Ȟ�s;jNr^Hs��F͍�,剴xW���[r�Z;�Pe�<D��?���< J���&�TL0;�p �
�q�2"�G-L�~Ł�ت�RQ4OX�:�ӬF�O�Ρ���[�d��G�IP���K6L&��}���p��;NU��6^�AS��t��p��B�?M\缀J�㭲��tO9�*N<89Q��\~~�F�=�7�p��V&�O�<���:Mגm�Dj��Mf�L�����'�gQA�-~���&&�:���>P-?�ϵ�g�EZ�A�xW�f�[��?�l�g*-8�(��p����D04�v����Ȩ���5ޯ�!7�	�.'�\h#�)M= ��J�NJ�iI@Ƥ8 �S:��K���Z-(�	.�&Z���^��X(z��R2o�t�����R�>�΍s�����j��c�����D�yC��t(�d�uۖ�<��㢲���x��*�f�P���`���be�b�As�A8�݂�f^?��Z�|q�k%��?Z[���MU���W���b���W�y�Z�+vs�5שkw�77�z�*�=W�M����3�h/�?��}n�v=��ț�	1�aWI^��{D��h+M�^���*4��JU�8�)C�{�N��1��1�x�;����P5L9�^ӄ��nP~Ґc�D�L����*pLUʓ�ۄ�ȵ)h�Lzr���]^�o�ڬ����蘩��0bFF��69�Q2Ys�1���Аs��
�J��k���5��;�Y�c��ۍ[By7[F"�c�r���N��RN\D��F�� �|�(dum�q�	����;�	0������ʢ��gEJN�ىl��ͺ:XhH�ٔ�3��X w!�Zr}��!��-l���Cb2��x��p
S03�&#�����O2��%����=9KG�~���l��/��'A]r4(Oj�Q;����Ȁ��&l�M���)v����B����)��ar�
1�Z�R�����dA�)��f����������e���3�z��b��N�{��	�C�\�k/��r/i6���M�E��㋢_/̻+R��wMM�x���h���*?iud�̆�bM�����[�5{<����U��@��?ޠK�p�Gs]}��"�[�u���1�U�!E��m�L���;�l�^7���R����)WS��� Л�g�n;�8�Ā������aN)�0;��J���s���ZD�_e�?���N�o&�E��*$���	ӧ��"'�x�y����"��n%ql�d��KM�P��)�K18�˻t���\�q��tP��B��f^�8g�3z2��y���k�p�V�QI�7.���k��i �20f�<��xWs�����1�$�"2��V��+��H�&Î0�ŰV*�_Ե,�ùt��霦�Lf|UEфF�_^������$�������y�|Z�?�)F'#��#� i2�ɐg��7����h�!��j*� ��1
O�������n����L�Z������K�z`�`�0�"rV*i��%�x1vt���176���2�c�-�((3l�҄X�J5&wC�м���|*=�_ r��J1�&�������d�ߕ�&�dn�{Q�i��Z��3��>G%p�#��*��.#D�p�i:-�%���� #� �v�(�[�F�b\���Ry�/������;����Ԫ���&f;�+
��^�#��b��<E*�:+�fKm&�,�ۥ��1_�٪��"4hz�=�)�Z�����·��. b</2ɸ��7�sx=���0L�S����w瓑�k�'8���r�SmM/��Us��*�.�w�[�GCcn�D�8<LMsS�bߛ��r�2�ڎ��XZ�1�t��8������;t$Z���v�rD�-�O�o��K㘓h?�@�� `U`�wX_�qW.ݚ(�5����#�ᛇ牋&�>Q3��d�դ[�P@F����!@���"���M�@'Yq�Y�p�ѯB�8�Fw��>�-yE����)j�CG޸Xm%�#�׳h��3
Qٳ^h�	�#�@��Cl�����@U�9ᒔ�4,�d!5� ����q�*��$��8�TӭsB.'��5�Z�����Q��W���]!��`�M�|��p��U�er�/c*0���w��Wͬ'S�5��Y"b�0U�Z:Oؗ�R���v�� ��Ā7k�vk7�;D���#�e�[�T�kO�W�K M3𦦎֛El��WĴ���r�v�<~DRm�%�y��2[[�S�G��;��CS�0���]�N���/���,2P���-ĲV�c�����{�r昻�9���Ğ$S�ى����`�v���~*Xb
���m��L�o�rT"�o��� ��{����{�s���:�5$�v�7�04XsKe�̬�_����ΑK>�*^��6��k�ŕX��wL&k���x0vP���F�;G`^٨DT��7���}w(�j�7�u^��Y�"B�~�n�����o`�B^�Cl��3V)Yn��<K<��U����yǥ�S��e2��A�g`L�+��NF���_�=�6����F1�+���9oRҡ3��y������I�����@� �]�;y1zES�w��C%nH�J�W�>�d�PQ��`;a����»�Y_���ғ��9]I�n`0���Ϊk`� ��JC}�LV�!���1�v�{��(qR��il9�9$�be,��4��$]T�"�񞗲����pCb���D�x�>�Y��"�i���.����� c1@��j6�Nb��Us:��C�8zZK D���EA㮚�:~AS͂pS���0���d�S��vc�L0 
,�:stE��j*�����G�RNY�oK�� ���m?�=?�f�����C��a��]�I�7IK�謊b����r�zgs� ���	�V [������T�F�q`0�z����R9c3���b��w�s��J_=c��IG���:�(�UX�.J�%:��[E�c�n]���g-Z���4�����2B��H�c�(�5�c�꣰����L�����~���+���M���q,�Ɔ��[$����c5`ư[�sQP�Ϭ�6{鬰���X�u����.u6��a�q��|�H)�Z!�sH�8cuG!v(	�?t� ���g�{ѯI!��#�Gt��K���Co��]� &���0���2E��맚5k~ۗ��,��P�u��bZ�r��S��+-����$�Yˮ��Gy������i�DeM3��I?�}@9Jx��a�^V�/'�e���:�f[��sѠ�'���]_�za��H�ʒ���YG����t����@�rb��cs�}g�N�{���R��<�p���-͎褬Sy3�5Lkp��G��*���z5e��=$��8�n��g���>4������8�,.�#NI
��%��b��p��[Л� b^�~,<`�w�	�p-�N5dJP���A�Nӣ �ë୏=���LŬIa�������&4�=���:����/e�X���A��(,�B��;��ϲŭ��'�� �m�Z1X����cx�Z:�Ŧ��'�9M3���;\�����r_?Ɔs��-X�*wE��y�������Q�0��T�S$��1S����A\]���֋Ƹ�QxM���2�.��{�?�S��.Gl$J��
����Z��H1MBǞ\�uQ�3I��=C*��ƃ�!�0ln�uM�!/7�]4S'�h-gA|!�?����Z�΂}8�wڷ?� �5�i�gx
���_��1�5^B�B�Tߗg\�뷤��AC5��k���]�X�*��������Sb�2��
y��+�+䳀�Sn砀(G���W:��}S�B/�J�m,Yҭ��g��f{uߊ�\0젘��eU�R�ZA�/q�++�����Sxw$�����M��� ��3?~-f��5�&ֵ6*�N��!=�c����=��C��
��öu^D�T��y�ތ^n:��4��V������!m�,�-~�p"�p�G�a��V	�Ƣk	�7ABi~5�Swy�G����jt�\�RZ�F�f/��Οz��G�SLCC)��K�]�8f����Y�~�L$H䃠�YD���ˮd��Z�}@����qw�?�tn�i���� hL��J�����7����?6_z.��w��Ҙ=K����c��(���%�}������P؟:��v�y�Ǘ91�TRKmofr?C����_�}��i����t��>^:V��I2�Jy��%�P�'�V m?(O����$2[<Bŵs\��a�@|��g�{$|J>��B��+���&4q)��.p�v���g���"�����ﵻ�0o��RH�^6�e�Ma��-�P\�����dp0��Ar�F��	r�!�ړ��� ��=0<?����C��=�����/3�����?���?�R���;�,��c���j�.��1!�jW���Dˈ&Mt���
Zp���(V����os^Hp��&��Ux����t �}�w�G�����`CY(/�q�r_����?"4��:��Z�SQ!��eg`�&�	�e���s1���_+�ʨO�vב��pq����'���A����`�S	���2�".<��=���eq���;Q���߰�_�z/��Dd�5ۢ�!~�����_����|�N�I��
.My��|��m��/&�G$(�~Q�o�:��P�$��.|���.AɁ
?�͚���V_wl�L�0�kn�hh��?�D*�ı@E�ŉ��
2��Қj(8�3�hO��sj��ִH����<�&D�����n�� �]s�gČ;�$)��֗va�+����? ^i��{�x'w�IL�P�bM#��3���6/���n�4j[`�X����
ٖ��`m������]
�l�dC���[�D��`�Q�Q��gg(���O��R����S��+YN$��[y!�hlWl7���،֘��	��qQ#���ے�I���etLx]őnV+��Ev�mXy��Ӊ	C]~L�sג�i(2�>�����j�d��Ѭ�r8NJ���H�I�{�]Z!$��q*R�n��8𡳈䑂U�δ%H脴MP��ܔ ��F� ��s��@����x쿿I(�3�ҥSq�RM����Ϯ�jJd
h�a�!;=Ñx6��T�dF�ȼ��w��t�ô[k��ޞ�%�,����.�BTdY�6bYV�-Ї�\�lR�|��LB�b�R�Mj`�L����S�:�wV@�i՘'�w+��fy���w`ړ� 
�`���U��qع1�Ww��6�E�.�㈇M`?����+�aX6�9�	��(K��E���1�Hm���;�$��1ܽ�k���qE��ʴ�e�!j��=Tir:�U>�&��KbԮ7GNr5�U]��=�����=�`����~�?&�S�9��Ĩx��o^��{Z��K�ԟ~��6���i�M������\o�g�����>��m��X	[*�巄��(�#���~N!țMc�?d���Pd�a�1����m��L�!Q�M-�f���Fp���w���z�w��z��(%��@-S�R����Kb�t	��7nߣ���(u0�pX���̡A�3��M٥�e���D�k�J�*p��[oi��+�%7ɟ�
���Q(dF�2���vv5�d	���H�*�?�h��)�h6����tB�LasW�s<��yb����$j���,�E�[r@��7~�I0�@��6h�P}����s%Ml�29��-����\C@?�"��B`���f�v�}_ ��[��e��Nd������SH�i$v��f*���&W�ҿ�A^i�� ~(����7,ns�'�O�Re����J=��#Ga�����c�b\���2Ψ*�)���4���D@��d ���M��]��/�%��jֵ�%�;Y����\q�2�xz����b8�v468t}�>�	��M��KL�6�-ڸ^T=��"�6��6S�D�T^S� ��U�?p��	+!�֡��b֠�.�-��K��*�u��J�Kf2&�q�?��>Vs����G�_�´���e��K�|Ǿ�%�j��������>�S�oR/�浼]�����r8�0��~�~[�D��[�y��ǲ���4ܵYN&���4)c���G;�"�6�i�:>����,F�9J��w��4�ɒ�����T1�]�� <��DGq$�n$����o0���#���`u�a��O�Q_JZ7~�8y��]��IKO�*q)�碮ڎ���d��"-Y^�m�	� zXgW�5ZW$_���8�ϰ*8{x����$�]1���ΐۄo���ս�C���V�.��rj��l�>S��;�� �h C�R��?esk~[�)��|����};��#}T��ɲ�I��9~����A�s/�k����u�"$�M�pV��k f�>��&�p��q����Q�z���;��-��p5?���4����RD���.��_%��J*�+e��c�J�;���I��d#�_�
#WD6�0�~ �c����i�iy�z6���m䴚!	Bx��Q\y��K��f��H��w����9�) 8l�
׈։��Be��o�Gj��-Ny�2����٬���y����`����O:	)�'�,���6m�T}RU�@��Tkb���f�ʤGU�W�"�O�$kU��z-�\������*Ň��
���/)jl}��yXy28��M��{����I���A�G9o.�׿m	f?{�n��mәu9��7�9�.oʛ.�����s�&-�Q�Q����n��Gu� ��QU�?u>Wޮ�X�#�x�Е	0��A�	X���-�9�<t�w��� ����|��+T��to������8��2yQӣ3��t�-�O��g@%F�Rk��>����k�ք������4x�د��~1%U�T�}�5�`�#���<E�n^5��t��sd�(��EU����r����0e�Y����0@>`"�!���S�L����74����0��.�I�:�K]:�ƈ5>V���:X��e��X�8;o~��s�  $o��3�"�)��#z�)!s����δX���:��}>�y�����<B��M ��O�
�~ݸ�Dȝl�H	_�����ȷQ�����h���U�g��b4K2O��9k�Lx[
)�;�1>���'&�6Rׅy�yz�&w8�axL��30�i&zߓ�T%��7KK��[S%��5�P����) +�˛�`iӅ`����H��-�X7����N�Xu��F�
,_��m\>z��{^Z����	�H�,��"w��|=�(U\t�rV��?�]羛��z�b��q�2��e߅"�[#;!��1%�D�1�/��؀v�N�,1L"{��b�s��'3K��ݛ��TH5ư|��w�����+5-ՉT�f��9.����pM~���"ӑ�7�}S��ⱛ��<�5hR7�1�q�`��2�� ���z�'��feW���_g�h�A��1hU����%QP]�`�c<u8��P�)�^�Q*t��+e�h.=ʪL2����om+eK�A��;p�h�ū����P}����sنY�r��}��ɋ?2`��KK��_B7\ԫˣf��SҴ�Zq\i������6��Mwi�ͦSڸ���:��uS%��T�╝�xJQ��?;I��y:	�&��u��C� ��`$�b�%b]S?�0#��ž�B�p9l�� �`�Q���[���v"���c�X`�G�k��y�����̀���F���sA+4��_];MK_��g�q��z�ͮ��w��R�0Z�'�২�N�l'p���/9��d9�c����]����1�^�X�<��K��c�,��jܼ�Z������Ȝ��v�G�Z6@9k��d���@���E'%L�E�]Hj�.t���
2��!��Z�r�h�����V�^��m��~Iq��Okƞ��@������3bo5�g0V?s�9�b��Ji��f������M�yC�v%��A�܁^둇6��P&�)]ꋂ�k[Wv���t�f%���.�K��]����k�3��&�:[��
�m�B"灍��3��.=�VQ���P뾱������{g��w(����]�j��V��81Z���O��Z)��O�${�^�	�����D��ÉC_�����!���)��{o4���QɃ����xD{@�#H�1�J�3`=w�`�FB�z��I��&"�v3��5=!6�����_��'"�;��60�bh��S���q���"��9�(�eAOG�w�U3]2�&L�l��
�!�/�Kx#�x�{�Л)���f��s�]�g�{ *���aϧ;{3�6T�%�|)p�6u˶ �@��t��v?��7�xs&9���j�0�s�8bkb7�(��-�"���x��+���Qp%��M?ּ�_�Q�D�:�"k�>=����nXI݁�Gb|�<���/�ؐ��آa���(ǀ�m6���Q��\=�=��Pz|�	�Y�R��xw
'�>��E(c�ݸ�P���Iǫ�*��u\�4J��ғ�ԯ�u��YG�FZ���j��?��MY�fs���[_���	U�eW��Mj��}�O=�����C`���\�U��&���|��w���=z}�	�v��Z��h��X��er3LS^?��E�����&]#�FN"(����6���7pG�*iF��n��Ǣ�>�Yy� �Y�W�Za	��9dt��@(y��0�,�\���R��w��4�a��ǘ�)ǅ|�<�#��ŨY�b>V�BH��q�q&��5�����%B
}��J��Rؑ���ubR&qT�0N�c�nX5k����TSS;��5���G�m��u���5�Y҃ԏ��.P���P�{��5\�����Y}*ؔ�	cI����E��`,M����a�,��=Rk�x�e0�����7f�����t�/��n�3�~��)p^����f�B�}*�h��e1�h$
�P�ݦC��=���iN�E0��/�R�f{�dlZ�Y�y�H�a�]�Z*���~���o��x	z''��.���`Tp��o�~w:��=)Q]��rX������q�n��:r��<�蟛@�Af��յ�xYh�M� �O��V>1n.�W@�l�}B���W_�J}��|F�/�/�$�K����6�Oo���<)?:ᡍ�uX���_}�8�N ��r���w�ha�\��V}�g����x��|��j��}J��V�ba��7���l�gn:"5�5)��g�%�T5E�k�ü�D����Lڡ��y2�����@�D��Y��W�V<�ٺ|l�Q2�� �7s�?v2��I*_������|�����N�&�����;��������<�?�["�/�|��B�Ѐ,3������ݎ6C��N�[Skף6�F6�/�b����F��+�W�Ы�?���>�CK���g�7���|zۀ��H%��P�ͧi:N^��	da�q����U�`��v>�$��`[��:��8n����;�5I.����~8�J&v�V�����l e����ԒI����8KD�k�������%�$r�{�t۲���[�=*zV|�����Nl��=ͬ�D��s�Ԥ�[��
I���ѹK���~c�9 b��ϭ��yz+���X"�qB�I�r�?����~�)�ɬ0�o�O�d��c�=��~��A�,$�	��^��
&��W�����?��3�"k� �D��m��}�����|%��۱�Y���Gm^\_H�������@ ��{/s�J��	�|o�;���[���6P��)�ZuhN}�2�'����(ػAѮ|)����M���Ĝ�<��
v}+�¢\z{��m���~�H�d���N`���>���1�E���Y�)�\�֐؁6���6�743$^���=G��{��S�A��(�c�u��ioЩ��MN�v�P��ؖZ�~ҊO��Ҧy�=�	�zS����XҴ���'�I�՝4ɣ�Y,������3D�
�YH�:�	k�k׵T6`e�I!��^�%�oF�a5�-O�k�d��Ll�Q_�`(
��ۿ@M~eA�L��R(�
yA����w�'�G�S����, ��^�EMIz.Z�����?�����D���f��|8���E)�F�$Q��)W������^��Xt����^��s��x`*n����cFb���������!� �e3*Č�}^eT�Ɔ�~���~@A���[��2y�]/A���i�����1���s��y3�&%����*B$_���@L�a0pK�=���T�+��*�L��G�2���B���k���;��I���1�P�M�K����`�G����l�ue��4������~/P�j_R�1>��e��*��L]~�<:��0��&�`��83��}j�ʚ�Do���+�&��|Sc���>jU����`VZ5��A�7R�Ӡ��>����`H���}Ӌ�G���D�%�?���6C�7��>��]������xT���e���u�T�Qۊ�g��1��'Ho�l�~�Wk畃�H>��[��2�%!j��xX9����1�(v�ۙ'ቶ'_�9����(H�ͯ�K��'D����]\�|;��e��F��l�d�1
{MF-g��UȦ��� ��cH岞m�{� ���o�vaor�9N�����vxĺ�@���zw�ȿK����{�b*V*�.��htf)�����W��ҝT�9Qo���6�s`���7�S��#Y�d�LlC��?@po�UvZ�-�g�Y�̞/�����q-�!o-�a݉������B�޿k��L��C�HJ�ޞa���]��5�.��zlvv�{+�m�X����˭1�!ź^���*��RM���n�+=E��JT��p�˦���s��A�BX��i���P�,�u��~�I�N�Apb�f��Bz٬P�4�m�p5N9|Qu�F�k����_A��Qs�킫����V�9A��W��|Xd3�4���>
y�D�c���-.���"D�6�*K��i6��uڻm����*�.��Z�Y�X���ld�/G�X�ǂ�u+@�HU�?6��1�^j�([i|s�V�Y!�����6q����ϏX�9�����о�Lv�(��!�}��,�	�.5RM�|XG�j���7�h�6�����h#��w�gꊏ�7'�����je�����eZ��[�aڦ�E*����{KS��d|9e�qT��ct?�j�u1���M�j,�	}C]"��	D�T-"{f�?�������{���5��&�6��=�ա#���% ����.�lWs�g�%(�xՂ}��W��W�yS��Eb�rXK��n͐iId���O)ԍ���$�UG�>jJd0�ss�	����]8mGwr`�n7��7_qarŉpZ�t�]����z�]�'y�W%�4�3*�?���Aeź�NNV�Y�fhpB����	��Z(�!��6t5Z��Ɩ�ˤS؍:7sS�pK�ʶ��b���	�Kpо�F2�2��D��y}��&��H�Z�ZL%m���w���[�G;<���.�5j����"<O:��/ ����ϑM�T�-��v��VW��Z���^�b���"��9QX��T	����U5�J�w���{�$;���0�
ˌp��Ʉ�!N���)����|z)P�Y�7��O�^)���sKx<���u6 �"�5Рg��>dEAM���p�����ty>�L5��6���Oi�E1�Lb8�aɄp�%���O����w�;�u;	�󫁥esWR}�9�@���԰
�O�����q�>�׋�ZMi�e�t�Cz-�R�V��Dqc	6�Y��hXI����y���(N�d�<������	V��)���M�P��)(σ���G���N8<[����9X����n��\&�9���6w�������z���5���d������R��!�:�E-fP^�H��	��@�P1#^�鲻����)9����L0W���d~��0qyB�t#�
�yMl��<]@�NJ⥂I�V0G��mVg�]iR�V��]\EWL�&
� �U�h�f��ЌI�3c��7V�/� k;��w�nI8( �@��k��E��8/���}��!�H^e����C\S-k���{<;��p��u�<N�]�/� �(��L��Ƒ���W��߈Q=o�`Ś"�3!`�|��C]��X/�I?��E?�U�-�Hָ[!����L,����{k��;2�ӚG<���*��,����Z�p���?@s0/k����L�ěUB��[mo���x����Ԉn�(*�+�z%�U(��@�!��a�����2�Pʝ�[�ak�	���g-f�c�zL�M���P���3��^]��x���:��6V�{1���UD=�����V>����ZL��.%��@."dU����*$���#���b�k���.��r#��J�C��?S]K�gikus��`���H�A-q�_(Y�6�[���� z0R�0��=rB|YR��gWU���4�^U�!��������Jw�����h7����ɝ�mzڐ�!���%�:JDjv�(=�F� ��DtP֊Zi��:a�Z�զ^{p���ˉk	Lm�L	��o�T	%��#5��~�Eq�� z���m���\��� Ņ7ݓR�69>��5=�gS3�����4/�w�� �����0��lN`ڄ�>*_��9]��oT�����rk�_`Ȅ��>�w����~�I�Y�eU(�S�~��-ڂ�!��q�t�HG��i��j}��4 ���|vM�`�G�3�u�;�,�5|��m\ȈV��.�4'�EG��1r#���ʵ@�R���"�9�j}.Ḅ��4�<&Q�8��߳�{��eԓ�����������m��X�g
i@j�e���d��EϞ(��Y8yFFǰz��&���<B�/���Zo�d�kU�*�
=\B���
�b�����������w՚t���\��iѱ���+��-Tbu[6��]��ڙ��yZ���jt�SEM}�SPو���։t�Sh�آB�w'p#�-B��MI�Q����a&�l����b�L��SOí�3cw���[����ŔB�ۃpGڙ ���<�~����;6�U���3��Z��ӫO���%���8q��H������)���4w-��4��)`pj���1喒�p��R;�/?c�g��yY[�v�c��V�}����N}�9������0Dnt&���t!p�����s|����z��N�۳�bl�n.B6QF���G�r�����CBz��ǘe[i\��m���l3��T�=��SK��7�+/L &�a*�sg��`޶i�_��}^��괡�ciֽ�5�eq �G��AB�g��$� � ,����udU����
D����?��r_���[�熵s�3|�mٺ7�KS���`��c�{���m�O�m
xE"�����'�|ye &����(��LŔ��3�.`�M�ٲ�[�t��`���8�3W�֪Y1$� 	�V���;Ԗ6��
��ڗ�b\�.eͅ�V�0��T�\LL,�N�|^��M�Z���&(�kj�����y}$�'��zU�&њ�4�@<������C�%��O�b���2{f3�Ż�fTI��{�)X�,X�I�Hvs=��W��s
v$楸;P�3�����f�cW��6J���1��?nˠ�4�A�J��%a����k�"O�^,�݃q{-�:�S\�C�no����9}��e�S��c�Չ������.�����?�ݷrS�
��LK��P �`�+�B��o���6��{_��=ѕc׀�dո4=�r<á�It�9�%:.H��/(�C�*D���]|Y��/�W��[���$:��^N�	W9Q;��hOQ(��^<-`��Hѻ%A�M�}������1��9��p9kG�K`���j��he�ސ0�x��@���
�\����F܈}W�r��ڈ�䑹U��)�p�a�bU����&Eux�Z��Qޱ{t"g�^��E?R��Y�9�����su��'w�,� O��[/#E����]%/	��Y�J!
�<i�1��K��+�(����Z��ˀ�p�>n j� �0�Ǖ�� �T�:n��9D�<)�c�����A�XE,!pw���U˱���&T�~�+QZF�ǄV��b'6i��[[q�P��񪱞�%K��%U�v�:�sb�� 2I ��n0��*�.�����}��q�ѩ��[�C��Ė&V��ф0��էp�L T�DP&"Mu��s���q;���Ĉ�/i�9�׶)��'kS��j9��{�7b��?�K�{���[_��n�;����xRH5#�IB���E;���\���@Ak�<�h���IG~����:��0]�K����Uk��
�@���Un
�e�|�^ ���?s+Ǐi-�[ς�;�[Ş���n�|�[M��!����[����M��:w�)e2��%\�����VSC��h3F��&�覬����7����-)�' t7F�;�<HV��
�W�A�8�r 1���3���":�o����ΏD�;	YJ����tR���@�aCOs��TwοY+���	f�Ě�=��E�������Hj3y�I�K��H����ނ�Cɦ�/��r"�i, �Z���@���C`H���u�;i0��o�|e���͊�M�=�2���k�"��mdx�Ɠ��0�SR�#��(}Q�e?�uE>�@o��^զ�Q<%�y����b�"*����a��,�STǡy�Ne
Z��X�������f��ϋ&u�x@P�/�T�ψq�����a�{����(��mհV���Z�8ƸR[���}�GG�8�	�U9�8@(������V�����l|n ��c�<$�y�Z���f�5�z�Ǔr̳�8g�����' �|S/~��^��.�nć}*HR~�����幜�R�� �f���(���V+�H�u"%b�s,��X���l��&��w4��	����� uZ��˫���F�\�����t��̕<��R����y��ȭy�Ʃ� �0'�����Ȣ<���{Ā�6���7M1,��a(`+�]r���v��c��*`�J����~���E�飗h���J����3�ȅ1:[��e�{��7����^�p����p���1o����j����#iE:�z��~�����Oٖ��s���t�"=䫅���)�5�����F-�{|�Q��7���#���V{`]I�h��kM"J�`���l4C�u����km�  �y����03���6��N >�����9���������s/$��y�f�ST���F�97j=0W�9f;���6�>cv^tNS��%�Y���D ]K뫆T�#)��WIu�yN��j��r����s�!�����]����.�I9��qI��*
�߽/WeR�'g�3�d��4��E����7*$	SqEp�/[S�^N��H�����^ܲ��u��E���eF��م!�*��v��Y�U~�)J��wK��c���N��U��&i���8:b��
��қ>�8���0X&�j���ڹE ���'��+5ر��HRF��Q,��%m���>-z����|�]��+�{��VI?�� ~A�N~��aQ�k���J��b� C����߷o&<��Zϝ�s6���{�&~=�ʙ�K����i1�Ʈ�A����D����ӂ�Q�)Ӫ�5o�i�DX_�~S���g;M���^�:@(���[ڊ>�ޘ�a���;����^���o��ؼ�� c����@
~�b�=0�dP4:���Ɋ��y�jĞ�#J�l�s2U�I�d!Y1��������\`y�N4e��G��:RbPo���uҠ�n�e�A�Yr�A`�5�K�mxL��܍s���[?����l��X�C� ��ҕ�-�����{��C{�w���`� ��d�X�|Asn�'�.i4VK��yg������1u�欐�����d�P�7[L=���?Ñ
G6�_O��%P|������N�T�<&7� �W�z4u�Ƹ�X�$��_�4�.r�Q��^����Nt����n�	��ל�T�`��h o6'�P�>T�a�I]�L�U��&2ߒ��v��T�"�*>@/�~����9��̘��<�3����a�<� �����ž�z�+臔�xP�b8 	4��C���4w����תE��$`I�(.�տN�i���j�EW��C&L��mU��l�����&�i �s壕��������E�v�CM�WX�p`���o�1����Օ�+@���<K��
=.��߲}o]�z8	�C�I&�\͠ t���ư�<Bˀ�D�/|H#Z�����T)�"|�v
���O�S��7T�m����Y�W	��v��yu��!E)�>��^ݶ�[ꡉ�k|��P�����NA�Ȝ9��f��q�0��w�+�W"� ��dD��J��<�euK� �嬸ξ����eF�������9C�хu�˕P�ܬ?H�gBn��/����p�ԯ����" R��V�6$�)d�$��N�Ć.��e6�ξo����hY�Wع�4t�|���T��U&���<�G����AX��u>�	f[��  ��h)�/c�C�za 3�Y54�PA��"�������	'��n�c��'0z��6�V*uW
����I�:`^��O���jqH�(v���\������Z�{b��q���su�@ǀ4́_�@��o��1�t=/������UB��z:�(Rz1���|՚4.}��nej����F�����L��e2�C߃S0_5�;�"�L�1*�)����e���vh�s,��r�=�Msm+]=���`	���ĕ����4CDIm���.�F:�zH�QQ�m�4s��ٷ�;U������7(e�a��sU���lޑ����mk(�_e=���V�mq�f�z������à�B=���m&ƣ��!��l�D�A�ڟ�Ȗf
%u`\� �T�2@d��#`j3�]#��c�&������OGi�mM���4)�~�}��y��qT��YƸcHo*�f3d>�,{w%D�ԧjykF�ndfq�\��Y]��b)��63�^Ӂ�#��?е�����rn��Cݒ�ViUL���&e@����� 3�5áX=W�"�J��{�q�&7�L����y�n�g�!��LA���Wt����,���$�+89�Ǖ��S���̄_x��cv�vE<TS��ц���?B����
��&���1�U��X-�����(��#��_�"�%��B�j���0�?S�Vg�[V�v�%(�fق$[w����G�G��v�O��Iz%����2��!���O�ʳ�k=�i-0�V�U��~��R��*�B���9Lj��%�!�dCb�dS��bm��*L��%`rfI3�7���Meί'#hȯB�8�z�L����~#�6��4�?���&�U��;Ҥ�$��z��)�4]���p��<���/bNTU�!�,��E:T���������;�� ��8�bu<�2}��v�x�"���g�>���l�ը�g���Za`����#�T����K�c�x�Y)�|�Pb����ރ�n�
D�-(i<zbSq����e�1�2�}�"�C%FZB^-Z�b=�������R�יr'��3��{`˨_-?A��B�x�Z+z9Gݚ��Щ�����a|�u���xjZ�"�Gh4"">m"��ߩ	|��lY�j��}��"������[����e��p���s�$���� f�����~�-3����qu�B���Q��&`���rW�6��o����?meZ�GH*cG���x_f�PE��#�WU?zm/c��`��}���8�:}Ļ��z��6]�q[S+��xk�7�B3T�@���_-JC>��oN�OGH��� ��6�G�2���	IZ�*�`q��A'�C�wߜ3�Y�Z��V�"�/`Os�n���G�<ߐ���>g�c�wX�C��5(�'M�k�\� ���o`v|��ZZ*�4�W3�lPvy A�5�c���Q�����i��Ѐ��k���C1��>@lՕ9�x狨�7
i��+�"f=kF���81����^�$ּ#����:��!���\�ڿ#)c�A�����=�nĢ�Z��K�Z���~���,\mX�[�>�9��$d��$�L�����(��D�X�Rp��%zk�*蒙p=M��-�����8>���	5�ʅo��.�N��a$�ȱ+E��
��i8���4W��E�T����}�i�j�<g��Xƭz2�U�0l�)7�P���C�ڦ���K ��XȡD�Y�g�S>͢�f�J{\ ?��8��]|�L/�J�;�3Mwa���=�f��1��e���-�bҪ��[��J�-�tK�x���i>Z�?`T]1�d	9�˰|�`%��i��:�i���)�ʁ�%ڰ��q����rЦ4��+��đ��e
�P��<�谋UX.�x��䄻� B|Q9�n-vw5�H1��(�h�M۷�p���*�Q�����18��y�B���/;(��ZuP�P+:q	��tF��b�>�1b�t��|[5�����k�NG~]��z��Z��
٩��*d4����U_D0JYT��g�莱�,���*̧`��N\��e��"��_�K ��4�}�I
��d��u�S+� #j��5�}q�\�U�D袆��
K8��P ��$gK�[�g`Ed�>���������XH��x�W�`�V���VGAz|%6P��;7��ڈ"N���]fB��R��AՖ���7u�ɪ�t���}�,����a q��=����|�� #��#���U$o**�{�i�3���D�����#Ó�E�K C�T��z舀˅��wg+ٚF�jO$�N��p�f��j!�$Ul@VF������b@u�7\��ǃc�9� �4������ζ[0�b�qd����MӀ��W\����"�3�i
��e��Vw,�4���å�i���d= �7�w��-%x�2�S+�[�nlw�_����9����������W�t&��	���h%P��6^0z��g�9�8:D��&o���?��g,v���.q���GoaQ�%v���74����VapASs��Q�3ڹݩC�X�x 2V��&X[���J+9����)�B��Z���#s��f���1��m��0�Y~����_� ъ�I��h]%*�P<If��^ݵ�f��xg5�6;�O����W�e*�#Sј�a�[o��{�KR�cpG�+���d/��\x��y���ܲ�u'�yO�k�����0��Y�&�C��u��ט�}nM����6se���H�h��#��,�O�L�U���[��Gd��rVH�'���]�}G@��-�߼���{�	��ҔZ�5l`k'���#=o{Sҭ�����[=��+��&ڍ#F���	rS�9[
�j[��5#����]EI
��nI�o<Pz���������I�;ƞ���d��ڮ��4�� O3�݄ÊŘ���4ן�-kWϾ��t�:"Fil�� J&D��.��ʓ�F=�?xj½>�9C��](����Ȑ���<��$iv�q����
e1��ì���*�0����������̆��fS��Fe����j	�+�ːu��?^�&��)�S�HXo�x,?Wjq������~灩�z(W[=
[����p0�����%1�������@�!n���q�fpc+Ы��*W�qC��2���"Z�� 1K��!�����6�v���໬�]��,q�M��g[��{�0~v�E��[���a�������s`�!����`D���.#]��_BB+�1s����(�)������v�BU�
an��3��qWA��8��<��(�?������~��ʆ!���!o�Kt��o�ۋ�Z�A*�k�F�K�U��8rE�?x��`?��� \��K�9p�xsFrxו(Ȓ:���g��S�-/B`5�Lf���n>�*I^�E���MX��2c��+&�t�r)�G�4e������0L���z\~�&j�����V����}b�l�]Σ a�z�ʃ���:6��rf,��~�;�mY󾶍��Y��D�1��ܨw����k�+���;R1v�ʲt	���m�j?�N�PSnp���G\4�+G;��ɭ%�,�SW"�yKe���ٛ�É�'�Nlj��ӟ��KmjHF��/����u��0�ul$��bZ<����تuz��xr�jG|�ݻ��r��C�y�˙�c'�;s1mG���PV G����wNy�+L`�o|��+�k�ɺ�έ��������P��.6���T����v_�tCy�L��CZ�����I���D���(*�1�
K���1��i�4/�]����7	�W������{�*���j�c�̣�(@�=$�/Q�-H�����{rP-�K} ����ܢc�S�b��,�n��9U���`.ρh!�1ɈVsv�Ͷ�R�a�	��ʳ�)(м���p�}��,�	�>FQ�i��ٙ�X�'�?���mHl����$أ��߇�a$����^�ީ]is� ����ā-1�jhY�(=��l��N��\᫴��a�wDˉ�歙76fDK�򱾥PU�q!��~Dc��/�ߵ�߾N�i	!�� �yX-<���D���vT����jVCuť�L	�^�.I`hSЈ���D��T>4�J�f����k�˟�M�>[�ab�մ�1��k#ß�ɘ��Ő�x�L��t\�=���S5�xF��ClV�cr$��T� 9]����R4`�D���x�a�_"��r��}����8~��̌v6��Z;�HC�ˏ)A����*���$J��˚q�I��ᑺ���e}�UT�Gz��5�Hu���3�L�,�����8:�T1'`�z2~k8��~t��O`(��� z���l_��r��P)���o���Ғ�Û�
�� ){�x��W��H�K �`P���N�� ^csV��+/^lQ��B����P��iۺ�x���#i��X�d`R���'�W/gR�yP�s�w��/�D�0O-�������Ykt>͞�1�d�>m�H�0J�;)����E��~�sow��d��,��ߺ^$S+�^�� ߥ�d�����Ηc�7646^�͐&2�z��×XL�"����r4� ��HϾ����ֱ���>q~=.4o�Cn/�V?�����|�W���qv�/
���'(�ƫ������Jk9������DX�kD�9'AdsQO8���'(����	��C��X�;-h�����7��G�b�$��H�;�s2� �?����_J麿��>I�}�۝ ��
zZ$8T�Xt��I��
Das\zP�/hJ۴�ê�e3�ҏ)���,�CWqX%�40�Uھ����p��u����������2Uz�+=��}s�߁�	�f7W���.>�b	�^�$��e*�s����2Ѯ>��钧���߾�Ja���{c��NC�ư���%�E��r~FJ�r����
�m���G��c�J��7�UBg�0�����LO�Ď�X�H��F�Y���	�8��31E<{.��.��{��$�X���:�g�[(\���M��m�.V��כ[��N�~�	�HFzn��`�4�-/����`V�@b��/�;��	M�S��B�MJ�|v����;jM;�[UhJ��).�<�S=�Y��?�vH�ms���7���,��-3W�v�b$�K%�e�a���#D�B����9u���X�/���Q�]��)��I�d�֔pF��|��ܪ_f0|����Zy�#~���_�D��c�`�^FlsС}�u!��͖��*"z �Z�x`qF �w���
��~���r�[W��.7@����~��	�Ջ /x�ǩ9�_@�r��c��=�V�5�y�KO}�G�R�c�BhOE�_�5��s���,Wq\J� �����x{�= _�T���ۊ�؇�0�0bѬ2�7��i���-�>�䛐ӫ{�Í4��,�R���U�X�����0!�+���]�E�b�g���3OM�C�m���4�@�Ut�	��C�^����lc���@�R ��n�:Xu�B�+$NC�!�/h�M)m�\U�m\�ٜ����"�\+@�tG6Y�HӸ���b�i��-%Ick�ޡ$�{UMM�hh�ɽ6����ǡ �F�=l7��@����[�!���.��¹���0pn!T�c=�*�B�I#�ʗ�"�v6�FM����(k=�"��� ����W�Une��
�a��3w^�O��&ެ�]-;�@k/>�J��T7�m`��\o|��0���PGc1P�lS�w��'�C�������<��8G؝ZT�J�PN�>@X�7�k{2o������-�u���o{�Yz~3�\��^�b���#�]!	�"Q�"���Bv��c�5����B���g��/�+w;�oDg˪�]PI�6oS����u��,�wara�ƀ��'���.޷�@PYa��d�囎�GNb�%ɿ��ZL�U�D�]?d-a��;R�Ċ�#5R�u���A���y���ag����m�k*m�[��x?� G�#�t���e�7y�� (�DdIѢX�D��(e-g?%��^�]N���Cs�{�/(�Zo���ڇ�����p��b�.�m� ?>,��׳���zˇ����!��B��5��x���H@�x��1�暐08���{0���_<�xd�=��]��̽�^��p$�-y��SL�L|&���:d`�i-���;N˛_��Fi�UM���k�q����-�/=�I��P������ɛU��5�lIP��c�`�g,�
��N����K�-{�*�`'jgJ�ya�V-?�B�(B�͠�Ҹӻ����u�E�"W��)p�F����8xެ�����Gtp��h��ڛ�if���)�ӭtY;��0׌wuV�DĀ>���G�ʂU��
�ڭ��5�z����^�nhz���"�@���o J14�Ǔ��@z�te�������D�=���z��E=���Aҏ�oY>S����3Z�Dw��J��JX��T�����L`�!��N����_#6��ܢ�Wy���}*�rbKt�����4�1 `�^om�hWø�r 7Q����������k�F���#��|D�絩r���!�!ټ��%6)>�M}�7����(Ƶ��L�b��wKUэp�(V��Դjd�r�}�b6�2���\uN|����4_��}��:��>���s���_4�;��r��I�g1�n�!�(i��������������?T��eOu&- ��"�����w�|,�.-)�x�͉���I��f�1��������#/� ��uJ���}\�r&� c���8��[�[V�F��;~y�盹p� _����s	��œ�mP��}�;Z���܌u�cA���\E�Uz9���6�C�T-l��I>��2��¤c�Wl��;{sQB@;�[[�v��˫�( 圄l����1��/�o����I����asBu����.\Ό�&A�����4��2��LK���Y�<�q<7�0�0T�z��M��~c�i7�`%���$�4hM����4z����d��&���:�;zu��L�˹>Y�+,����9
��p���&�Lh�N`*#�����%#��,rn�*���Q��L�#��%��IA�M^�
 Heg��r�F'Q-[�[f��=�[:ܗ��ɭ���)և�1\9��6�&P�b��(:�ڲ3�8`��K8�/O�k�_6"�e��N
J}AF�0+|���3iۅ����)��h�'p�p>^gI������>3!C"��ï��Ϝ�6*X���5�7��ki?2o��.�l�	�
��f:XH��@��ͧ�~[恜�X[���%����0��BS ���,m�.Q��������Q�j0���n�I��@hG��#����أ���TmȖg@%�|�4g.iK����a��~'k�>��l�n��> �*�yKY6@$�*��Kn�qt>��{3��rܟ[�K�)��Z�����~�u+����AN��m�z��蜛!T+�}����C����y�`t����E[��(��淒u�4؁q@�,;�{SY��p�����Y�Cv�i�mH�����*@�o���mc��R�UQ
	5����(��i��y�����&�+�ʢD�-�B��	����	�0��.j�������O��th��AC���I5������Z��h�9GG�*�	��0�ɸ!}��"��<���C���hnNy(S�e��%��x1��~>��k$y�Pb�|n\#��v|��]ͯ�u�Z���������nX+�l�'�����(�i�l8�����Q��ƖG�����^mv-)�^��Kf�c���i�AA1��:;��� ��eH��xj�5/�R����q�wM�F���Ykŏ����{���	 :\s^�]�;:����)Nz�h
G.���d�D�~��G�~ ��ʓQX�}wv��R�8��d�;i�I�m�b��Q� �.]3���Ҭ$H���Y�s2�2'KC�k��Vs�c�7�*X&	Lvjj9���EÁAM��I�f�O�,����r$�	��-��v�|Q��q������U���&ݬt�Ѫ�z���ٓ�y3d<�"r�ItЍ$B7n1�Q�Z
0~,.�1�؝|�hø	�t�L�\�����/����-k_�,�9�e���%VI,[�"�Qh+�L"��O����K2�$D�E�	����>p��L��< �Y�R)�0����pU͌Ɉ����^@7���<܅ԞXQ���-i��Ѿ���\��W�nv3{�|6j�u���K�O��Y
�?H�o�S�jZ˖Z,?�� �i�2#3�8*� =K�e���s ��x�����t�=�8���	\}yqj|[��$�����߱�|�xmf�>i����#c���:8���=��n\��dتw�|��C�^l�$�k`5��^�P�cH8����"�<�W��kH�&�_��1�7����Mg:_6J#֖q�=w���Z��7Z"�#�7�
�񚭭g )���W��g8�A,}&S�R#� � �����~�=44R�C��ߘ��!��e,;���!��Ys��.�q�P���� ,�����Ld�hǩ�m\?��b�v�ԛY��\�s⣺��$�-�aή$����n�}�͖{1��'�)���#Ii|U.'�����A���
���:X9�K���s �G�d�	R�oL���NU����u|N����B"�ǧ�]eѹG���L��i6;Q�)D�����A��#�V�Ƞy��8��j%g�eQ�S̰�4j2�V!��Y�M��%�������3��Y���#� Si��$R�d �?�3�:u�)G$��I7}�~	���Ѐ�o/}��꾸P���pr?�9"�fEP�Q��)��^ԗO^��w�8+��\�HQ���ު����p�!�����~��LU��N0�:�Ԥf`i@��_R�c� +n3��Ϗ����򪷊��_a��7�K������� �׉נڇ�j��m@�_`�b��Ȑ��/8B��UHxD.�%�)��I1�W�#�T�$�ƅ�9�AKu���������>[��;��`U�}�
f<�f1�or��޻�	3� �C͂ڱE��D�Pn��Nĉ��T�����Mx�u�Z1(�i"�R�a����%m�
bkI���n�f�G=�H{��o|�Q8���唧�%�ا^���u+AQ٫Q+���+wF��rQ&�J]��R6��%+�yfT7H�d�����k�2�p�*�	(�>4���n87��Q�0TCG�cB�0�м'������x�o��K�;;�����?K���D��T]�Zx�0oS��V�(��� �OX�_�30ODO��N�z\�~�|9��A��$=��� :/��M�AQ�"ш�ŀ^ ����8�ad9��u�"FD�m�%#,�8����;�D�䖧��p)+��D��zDP!�������V�Eef�;�3�5���C5<ހ4/�K4<y�a��\dG�8��{�mL4��sBe�L����~��S�ߏ�T�ӵ�߁���UP	�Ӡ�A���X)�d.P%�Pt4�
@ ���B�|vfD���M��3u˓�=a\���G���>s4�Z�2mr���L�^�&�l�Z��	W(D��U�`4�)\�9���W\�8�����K���4L�^��t�B`���=�*��/�����{�M���J3v4|��cpJ[��[�
�?�:�d�S�"�����MG���g�c�kv��QL�=0 Q��̻88`#��k���B?,�Lj��9��Xi��-Ҭ�D,��Nw��FZ���q�)�H֫��ŗ�xZ�M>�8л�,��T�6����������$���>Eҥ-���g�܁��os4�VM� �%|�*�'aN��<M:������4cP1+�}��a^�d�f�	�(�����;�����O�U��/�|$ev�_l�z��:v�����T�\��<"(��>p����3=�q��4�c'a�*��sv�3��Δl �5E�[��0��>�oa�*��W��.�j`5l7Ŗ���>�'
���)'ܷ�rB	Q�T�p�w�e�Kj�t�ʯ���Ju��Z�i��BKP��,e��������l����G3�|�o�����F�Ϝ�7�q�%�I4��S����R�v���6d��zD�y���w��B&z��Ir�8���X� Ӈu��L</��>ȇ�ľ�M���5�p��o� fx�s��$C� 'd.����eJӡjJ}�S�ۨ��vy�N�CG��qh������1Y��:o^!�&PC ǷfZ���ZhK��X��MDq9����i/��-0��/}"hq̐tF8�lω��lf���Οy�ƺ4�X�����h��|2i���;E���F��Lg�Ls�'����ի��\����"03�O:�{3�TF-W��qCy`�/�[��)��H��B����֜�Qπ_��/w�=R�P��Ȉ� F[B�8���+��,&�/�c���#S!��l*�r�����)�G��0fғ8�dB�3��s���	�{i2��kp ���`űK��7�!@�橮H�{~�k����g��J���O		�&��P/��+ 	vyO�:3}�v� d1o����Li��#gO�M3C���s��#��-�������P�A)�6٭;�;�����w������2�/�N�A�c�h����nӪ��,�Sl7~[]ܥF(dtSJ�A���jD��ܰpH�ђ�+���Ȋ*������#��m�**`���!9��+��0b#�����+a7,Yޯ�!*��ގ.'O��`t�1��\`���:��?+����Zh�ф�T>��Rq�UGh�Pȿ��4nVV�Bzv�%Ve|�ax�/ԧ!�4�L ��sd-��j\:=x82��P���O��s <��H#^p�2�o�`>���f"�~���/B�ۦ����p��v
�^����&�[&b7��T����� 9un=�hju`�Y�����F��!�0�3>��� �;J��۠�:�~~@��wIͿ	YO�B��%���*H_���~�8�jD<�&&���f��hI��z"ܺ��><v˒(��mR��	aP(���]�)�ٍY��>;H$���@ڑ[򤘞� ��fA��iK�t�~��Ƞ>���g=�Ȱ!�w�q�:Ǧ�N��1�MO�I�K��K'$��[8�|��FE��F�$A�A@C�=�c �W���[E0�b�O��2J��	�6�90e*5���g�ꖮ�X郍�a�ƫ
�.ph����e,�zأ��͆����H��PCJ�,w/t��Y����?쌒_���L,���e�6������Ů�7B9m8������mN�����f��_�����U6tZ|���C�9������ҶT�^0BE(Ҋ,ҏ�$��@K
��p�}׳��4��N�u%���O?�X�k� b���?�;㡹��r�u0�:�@T�$�iT�����Ay�V�ޘz�B�����/c&q���I�/�D�<'���1_q-宮b�[z˪�H�tc�|�6�>�'7xL��B�m�c,iT��ԑ�,���JjUc�j���i��r��bJ��:�b�
	%oL��s��{��9�5+T�K��mɩX�_B?ew�������b�m}R����� �wIB���&8�V���$j��]����`�2�����pFkp�j�o��VB��7F狀Q���.�0�X@�7�w�"�F���d[���L5���36wE��2����ց!�V�>���8�ݝ4Y��ϼ�E�]z��)F��u�����L�U�Y�Z�"����D{3�t�퀊L;�8��ɓ��t�p�;ʑ��u��	����,�?����q6�����
p��/	��Y���3`G���v�)<�^��j�]��!R�`=�	�On\�<;>�E|݈d��w�a&a�N�;�2n�'���wx���5[��P���ʢ�sH]�RN�=5���:jEvNa�J�q�g�W�U"�H��8K��枸m��������''�5n��j87�셿;ڍ�H�2=�\H�2=��Ӗ��38�5'�5��$kը�c8k���8�V�:�]=�\�[��dG��
mP)��uC9(FIG����n�HJ�^�����I�;�l�#�65J���d���je7M��b�>���z�'��1�#�z6�.�l�ej~����Ɂ�g��	.��ȃ�ǟ[6�����Up�����~��e�v��eT�l�2&��iyW���%��lN�C.�&J��Y�.~V�� |
�3����kA�D��S�bp���.;Y��X�����TR������c�щ�7�c����f&I�L�\��a���2,%�����!�Q��8x��_h�L3����X���5�Bi������[�e3��ÎB�Ю�ޕB21;J$4@ͧG�m�,�#]��1#9*��#@@�"���D+��b�5��7���^�ѝ�Q��0�y[�P�{&�%t����Pn���q�
�/	.�~TݩH��Tľ�A��$}���Ώ�a,^��[�̑�_��a4Nj(���
���r��T�w�#H����W��Wf!�L�uC�b��(�f�H�$q��\�����1��:WZۜ=���[�h�#B��bN���`��j��:�����n���%�×gX:羋2 ��~Յ.%�6mK�����Cj���>�
Q�h\ua^����T��=>{�ڏƸU���>��^�‗�)��h��|w��b���Y��)��>���m�꽥p��@W�l����H���={��G�K����o5����K�k��1E
�E�W_��p{�0YU���#�Yߙ~�pWp(��� Ύ�ʀ�*�VòϾ�:��������7���卷�14Ʉ���N�G-O����n�fyż��u������x��mh ��@,v栗�h���0$��m���J�7W�Ϯ��Pꄿ �099��y<Bg"ֆ��H>�e(g�xLs�5^�P������.���M |g���U���ck�B�i4nq=�+t�pSK���3��g��Q����Mb9����Tr�C!A��c*���!>���S��d�ǐ ��&�> �k�{�����#P���O`�X?>[��5ܬid
/��[V-7{��h}�i��ǢΧH���
BmR�F���Pn��K��y�J�PpR	B��`��N8I
ӁsCI��(����C/�/S�ctP`i	μt��X����q�����g]aˀt�)Ϝe�E� �`<[F{8�eQ��w����򜰑�מ�7'՘m���U4���ݰ/m�_��	��	��gc[�j;бҬ�5�q�FKBϽ�1�Z;Oo.����ZҞSB��@���=��k��"�:�&5$_��^�f��j�I�̯&��c��>�{�y�T�UP��S�|4� �7���Y��VM6K�z>Z$�rҡ2���(D��h�E���W/�ʙ�*�xqqP�@-��9
��S��-����̰M����Q@I!~-��_N)$ɴe�ٿE���K�6]�S�~����v́�+����X�
3�~������q��-̶�y7�Ù>f`�1MŠF߹������=e^ϖ@���Z\ˋB�n��݃���� ��GwI���t�G�������&�C~�i�,J2J�	gש(�����+����ew3p$�2�G��:%�`���;!.`S
.Qo1���7��Xd^\�RR�6UƓ�ފ���E�G`�Jln�%�?w���4�m��i�c����&�1��9Պ�d�w�����S�00:�x�Y�l�7��k@Fn��MnW�%����b��U\���W6�EU!ܦ��ܕz���9��\b�/s�>\bEai:;�S%;�{������@�F{�=�?i�� �o��	!�bp�'��j�.�,�^P���H�1Ɛ$o��d&����EE;F�W�;c0Z����iݔZ���`�[����b���h)o��Gu�Ä�	8`���mUr�ǆج<���x��q�T��p1�|!��
^ĎI��Xfv�Om+�p�u�����ߍR�rcO���'_҂(����w�	?Vg�W{�)��X2�V��d�N"���&��я��i�y�0�O�h)�8���(�'�cG���z��o`7�a˓3�
B��,������1e�]�� C3�9�	�yH+⋁8/v�����3[��>&'<�ya�@-�f���u�.��h����8T	�D���{�1R�yg	a:�1�T�To�E����n��d̗�Iب�h=r���i�	;+���T��B�#n�D	�a��cr��:��� כ�A�����=~�zⱭ���x��F�� �rW	�OY���h7�".z��BM��J�h��4����1�ږ|@2����@�5�Ԟ*��))�5�SpN�z�v�c�3���S���GC����c�T�� ��7�ȸY��ޗQj)z�$݆�o�����z$�N�0p��͇,{g�¶wJN+�D4�6SY*-q�^4�v���x����އ��Ӧ��To:����2��{��$Eu��y*4�𧿀1��6�o��W����g�̈́y��4o���+(���7���)}kp��r!�x����kKcA]��rG�V�~�l�8�����:5q�_>�g$`�F�U0C^�˒>�l��f�#��0!�UW�\ �|'����v��@	h�C�3$G"\��)Mo4��������P'��?F��=iVy��B\{2��I�����C�ŴAsWD�(w��6�6���zU��������=���S1�Etyu��
��$��b�,�����'q�N����bKl<�E���yw��l��m�&��I32��	9@���a�c&z�� C[L�����v�7:0�P����G�FRRFp��0�iP_䨧�EZ(����d%������'�οM�ù�j@�r�;�r��>,��7/��7b��jyi�;b��Rp�y�1��w�zI�F��È�)MB6���
 K)s(:E����=@��B-w[�)=���L��[�
��\�ɨ��8�NmoF���F4֌ݒ���[��ڮ(�X�$	���5G�XH܏I�^���Ws��ב����U��`����׎V�Rs�x�}������R��:I��-��	Π�qo�u�����(0p{��{���<6ɓ�����_9�c�9r��w�W���]O�^R�?��t�D���\�E���	���v�"f.�K����W��x���[�dx4��vJ�6\x�Z���k�ѳb�
�ΗN�R�Ҫ�;&՘��{�_L���W�$��%�(�?�o���ｑ�+>�ȏ��bf�2P5���������� 
�uyN��уX��<4b!�� iɱh-`���΃����Z�b�g���aИ�ʏ�w�L�49:i�nn�cp��������p��&��ux�cy[&T����fG:h�~l~�4��*��f��g#.�$�J�kCϼ���6�̢���~�K��et��X�3�<�t�g<�v��V����=���q)Z��P�O~���;�)�� a��\�Β�N/����u���IS���i:�r��Q8�r�Ċ�'w���7���xq�b\Y��Y�0.�;g�{.�r颖7x���:�WI��U��N��/�m�j8㟋yb�N�劓hQRÕ�V!d��:��_`8{^�Z���\�*��D((L��@p�g�!�)k��F�����5�X�.�u��b (�ܭ�ء^a�~�P�_5�+ݰr�&,c�k"gҕz�x�3�ћ>��T�\i�"hN�)|
��P����Pۂ��ő�KϙS�J]�N@M�v+݀8�&��^nEܬ��r����W��U.�Z*��^wL�<�!�Լ�8q|%�|��HY�W_%��<kq|f�\lD$
��y(�%I�$���=m'`�:�ñ�2q��1��Ec�l���kD�WhP�(FҢ�d�Qa����`[��h<�<eQ<SI>g:���z���[��_fe�k�,y���2�]��/���5���Xr�Js��	��$�=��j�n�vH�"�Õe�X;�� R�I!�I��02q�6X�_I�޹_�d�7U����!e?+��mY<�)�����H�f�d�Pk)�D�H�nn���[��$��2#�a�>l��k��}��gsY�7=���ri�*��*�ֿ����/�L�j��eM�l�#��`�2��[����0��i�1�r�b��XS�%A�b�]_|(��A�$���Ѹ3����+a�Ax��
Lfiz@���L�T�b�N���P�R��������i5����
1T+?,�bB
�-����_�o�-H6p;������C̧����ngD��`)�L������Y�V��������nk:'_��Q�u��@/T{G�0)ߛ�dR��Z����3���ak�٢�[��jS����Q�Ro�+e'�3�$l��,���]L�S�֢KQ=��?���J �������m':��0���B��G�.�(�Ar14����z�
�=���M���8 �X�� ��s�1=N
�
m0�d��M]n=�$��fNtdO`�'Ц���Q&�K4��]�c��]/�_�M��W�x�F�M��U�{���){��O�Vw�9u��=@�<�m��J&Jj�@�� �(�!��#=��QP{�1%� dFf��Ms���\~�|������j��y���o���"(�P��~��,� k��@O̵z�������5��jyCɘe�\�5ln�����$��/�82�_��/�o�PDl��+(߼�+��~��{���/�D~-�O9S��JR��Of1�?��_�rˢ���f����Y�yÑ��3?��kA$8�m��%{$���q�8�6O�ܥ�D���}�I�e_~���M_�@�*��9�n�HƦb����"=[JP�;���]D�\,��t��8O��y�M�u���֜���}3�i8�~�'6-��L�����}�(��* ����ep�I�H&��u�0u���!6��;�(e�CQ�E����8O]���	&õ0�{�W AP���(cUvUB)]`�ݴ�7�7�ʹ�	mg��u
MR�%������'E���xj�{�J"�L�ԝK��&9�XCJ� ���I�Af�p����SI�"���{��uҘ��q�L���ef����k��@u����"۶}�|�
����jW���<E����1�����#�miQ��ȆƼj��q1]oz�T�AuRT{tN#��ڱ������ho�P����	Z��{D���J	�L�&o���P����\ީocmn҂���آB%Ub7��g���R&w�������kw�Ԇ��ɠ�M�z_Z>^&�2_�TMx h���������-��� ���Q
Kcߥ�H���x!�$�{$ θ[��U����M싇���N�[*��A(I5 ���|�v���=��U!C<f;���*��]O�d��s���br�����s! r��+!sZ.z�M/�����@Zx����p=��OZ�,��b&Qٱ73!
h��0P�2���������|C)f稕V�gY�4ټs��e~y����T���%I�Y��	<]D�V��ө��vuD���ի#�L]í�Y,帿y9H�`�Ey̒�kzc�;ӛ��S�q��隮�-�Yz�����(��8Ũ}'PU)�����9�7l��sTOi��,�*�lo�g��՛8}���z����'ȑC�tW��P���A�g��a�VC|け��r����h���~m�s$΂����cE� ��Ċ�W��}��h ������q��y�	#Zؚ�F��x���IY<���_^�I�oe��%#z�b
�G��М����xc�>���Ft�@�
�E�}��0�1�o����I5��8R�l:)����pjh^�����PP[���4���5���Y�#�~����6���H-!|��L�_>�o�Hm�0�8,6�٭�r�t�����e��7۞o�V4�ì��[ᯔi�߿G���4"ه�>�K:6������zK�s=��D3�9�c��Y�f�J���l�*hYS��q�1�z��$)T���Sc�X�#���hW�}�㔟�9*��h�����\�	g�E�b����:p��k--YUĹ���bH� 5���b8P��2�Y1���}j����j�Dp'I1�f�ޠ��(�5D���Bs���5�0�m�s�����CޜX�.JE��ԧ(��W�U_$�A��L�BD�c��u]ws�D;o]k�C�~�h�l����_�����<�W�%s�CMwS��7�v8Ћ����XIY���ى��μ�K�Zk��P�7�c���Y�)#��� ��h�&⯶֏Y[V��2M���g�[���)�J:)��7BJI"�A[O��z䇭�X��gW��N�@5��Y��w�����UH��d���<^���b���m!���v
�LQh�����Td����9� 9�"mS����D(,+l_s�HZo�'�?)zX!S3�~�'b���포��c��ő�F������^�E��K�x�s�v��}{��I����[˥��	Ї�;r��R܊�:�-�&KC�'8�Q3ZH���I��x ��v���i;�����؅�3@�򉶊��J��G))���a��<�)��D�J?u&���6z�jA�:p���4�kD���
�]E)�;�g��F5ͤ���#Wc"+i(�!m�i���Hf���rk���z�O��t�`��W�����Δ_|rF'N�P�6��� ��'�Y�����2����'5������L����l��sr[���x�eֵ*j����7>�ۨ�Xp�k�!'��x��N��_��*c�T�8����~cŷ��T�KL���� _���^����B� B&��/����ڸ d���S!��$��P���4���BX�6��!3�eXs�d\�G�S�h��Y���݁�o�S��͛�ѭ�͜�BW�A�D�C�ʺJ{D�G�r'RGD�
/H��/�i�,
��E��i�(�_����&k���G�Q�����0�hV\��:%t"��Y����`�Aj�3
�'r'��2n;X��4��nqeM�RJ'G��aT���^��}�L��ҁD����OI��9ڀ�#�>@��j�$v���d��^TD�&���I9-i�»C������3��o�˕�J���U�!�!)L*5݀u�	��6+�\�ax�X�`�HOa�]a���6���p$�L��F�S���"�wbQ���Iw�=m��5��DV�3~S�ce[��ha�����7tฅu��
��`|���7[�[*̼�c;R���t���xE� mr1��i&��b��ܢ� "����tg|�� �I��1g)v>��bz3��Z�ruQ��PL���ij	KV�W�[6�_
l���i�&�}c-�&�q5#�t9]$_�߷��CpyF�ie3��/���s�i���i=�XaGoI4�{8��e���ۂ���u�ʪ~�H�#KؼXM���Iv���x��-�,�Q�؁�(}obA�b�%#[&���v.�B�3|y�轚��M���<ȅ�XS:WV3.� A�^v�~��ɇ	{P\GȾ��	ў�v,�Z�Qlg��O\�n*�3L�
��dP�2�ZeO��p�j�X���@�Zk��U�(zu �#�7�f�|cc`e�g�0:�haDc(����0�_dx�M��l9b�s#7q0�8�y�{_��3�1����B��YA#����\��s�>Z�]���g	��ګ�|�_�bS�z�� �(�<$�x�}�#��v�z��Nb�@,_�G��8k���|�&���m��}��FC���f,)]����2�s��Y�Px�#wX�خk��K�k����Zn�5LC��L���[�S��lJ��H�v�޸�&޶f���Q���~Z�� B�ɥ�o/IRU)W��HO�cOY4W7ތ�9v8�%<�u	��]	���q�cV�f=�)��������)1
ȝ @�t��U�8��!�
$�gN��LN�	I����K��8i�K��W��)A�w42 ������/�~�-Fs<����%�g�)�,sL���s�\�i>N�;��\�YEB�r�{9����ԛ��۲��D�ʗ=ۀA؂.ٓ�'���U�6 w�>�y�2+�no�5�E�����5�\n&>��bǕo-��*[��c:�݆2�H?�ؐѫ.���!��L���5(����)t+\�14N��Jn�N�e���Bs�'�g��T>�8���8��'��ݞ�PAy�l2\���ؤ��j
���r
�P
�h>VQZ�c�PP7 �φ�d��7v���݊_b4����o{\v�چ�DO���~�h�1��p�Ţ�\#�����c���p�zT��jpq����V�W!@Q�ٯ��)0��;��r���R����J��w��T�N�"ndzq�a*�3,��w��/��1X��.띚����SΛ��K��#E�f�`4zM���T��Q�P�?�������2Y+��Ӝ\�8�z��0+*��A����؈��zt;���y�q���X�8��d���@]5�b�F��V�J������ �S]V�i�]%���2]��-�-3H�?�걈q���Ł�؈C����4@�� �C�kl�5������|�[s�oV���P�wu�	\�ÎHUA��9w�H�7S�? �P`��x�G��~��,�z%o�=Mf8o�0�ԓ�E��z�K��`6�0~Ü��X�du_G�8QH]�[�5����Vr7�&�V�>�,�[��B�Z�	e(�;�0-����Zc�)զK��ݑŐ�V�s� B޵�ւm��4�#�aC-��H�9q�9�oG��4��:�
[3t?"7�5;у�ӧ����X-f�]��d���w�k����WB����$�&ev�a���+5z'0�Y���V�c��+l#.�Á�k��m�����q���G#7[OKpjR<;���8U�`gP�x��&�N�3H�K}��Y֠]9��Q�eU��AƘu�S��Z�ה���:��΃�5u���u�O�����,��m��h�Q���+�u��3d
���8f�t?��5G
!}*`�����z��8˷3��͋�꿗��
.� ��m�9?/ةu�����5����'S��o2�oW�9��.��ӡ�5�E��[�Q��ҥW%��l�-�F��	''�������Kg!�`	�6�O�_��Yz�@� #Id�.N�L ��ӤX�Bp��5�w���n�nV���\�{����� "�N������@�$��*�y�^t�6�/���^g�?�ϑ3����[^�v�a�J�sK��^��_C��MV�J�������KF���?+���y�k{3����i$B7��!��Ț����R>!(�[=$p�X��^GՊ��B�S�Ւ�Ro�
�@������f��e���Rg�!_�h3G����>e�i�2��lCt��B��|^7��|�psK~_ޢP��)u�+�>p)�8(x��OI����Ǚ�i��Dh�<Z����Ww[U+c3�0���G2�Q�WDǭR��I�a�L��u;-�N*�C���4���ψ�/n͞�R����X�/�7%���5�۩��
�kD�Br����7;�.���&�;��o"BA��*���|U�2��v.V�Mn���$�{4ed%�/�d��5<�=r��D���]^���y�ԉ����mԍ�j�c�=L�Mc�B"���$6���o!E�}�(�Wq1��O>l��uǸ�����b��;I��/��:���;���|v�m�d�j"d�6�1�!��1��ԭ�|+�6�G�N�WKb�[���G�[��l�5�jGg�Ӆ�-*��T�BXV L�
��!�Y����u\�Ś�j�d���r�9j�%�0�U
j�;����~�6%�c���[���[�q�;�i���7A�y�!}����ϡT�����Q'꼸Ӳ�3%'U�וf�:�q�KD,��7Q�ԕ�x�I��-�i%���'1��CN�Uy����o�ot���I��D��z	-��}��]ʟ��H���{/�3��9f�
���J-o�����%2@{g9��ʗ���w�T�c�u�\��K#��G�
�6�G��r�gU��[m_9�[�ZC�(́@�ѢX�O�{hN�&;��ആ�p�/j ,}��� ��K\?~�*i~��_f>�/M��zBժ�S�u�T�R��,g�O�'Ǆ���$�K�sO� ��x�p��)�%9����a�5�I3�:L�Z<�CO������/`�v�24�B:����˻�d�a�p�*�B ���֙$&�GVBA�צN��Ӿ��K����(�=�rT��̘����e���=���e�x@r��7P��+��QJ��"7W���`d�W�]�WpWB��r��v�MW�[-�8�y�8�w�\Oa�Rp�~�F��l�#�W1���Y��P���}�q��Z3[��('Ǽ)��d\��kr���Z�=��ൺ�4��a!jP�Г� ������9�|���bH�,���D^��rs+P&�|I�-4L�������}p�LR�1`����R�.�w�֟R]~!��;�:њe�l��5�#��)?%������>��_���~�6��i����Y�rTȗ5 M��8��&���rf��)g�����9�u������|�l��K��"�w5Q��O��D+�Y���g��������$*��:�2h��+�z��v�JUGUG�rk��?��\��1�b�W���[���d��Hʚn"گ^7�ɠ���5��|`S�|;��]�YkT��3�^)�/��✦K�m U0�$�`���v��MD��U&�vt�E.�E�&F�� ��X�b D�bK8��� k���|�D�Z�ި	���%o�JDY��<����A�7�c���.�g<��&{����'��V�0�X�@<�u�Y\��K�^< �L!�`b��)>љ�����VJ�S�`.b���3�+x��,{�0���;`���nv��:5)����,I���?��i���K��y�ґ�Iƺ�G�n8�N7�*`�(�Mj�A7�%��5+�?�Į�,���'h��&^<|({EUh�^�9@^r���I_\A~Wh�/_:�������ږ=S/s�6�������T���h�6'(LPbg���
v�N���4�;C�6<����o����n�ZY�Z�J��Ct�/b���"*�<�>N �1d����A'�V�)���_������/�����)0�D	IC�l.���-p;�b�]V�Q�PBo�3�0��jX;��.���w~����O`Y;��X-�ֳ������U@]z�O�a��D���m���*��w�`�'V�m`#��|� Nͫ��� B;�<����FFg���U��w�ֱ�@7C���_�6hyػn�H�(s�`��{�R�Ԙ���[����$����㽸R�N*��4�1��W��ٮ��P�.Kp�\�`�0�K��k3g�S���;��U����2���N¹ h�&,��.m�nR� �-�/?۹�<��D��I���[Wn�%@�'�� ��y	8�6N+�YG�"h��a���@.SX��H,p��W��I!�6e���7�ڢ\���a|���/�ycp��7i������(���;GT	Ԇ"��2��J�답�K�I�tI��ȿ����}� F�����I�&d8@�uA�_J�)1�VϹ2�#M���EF����7�bԱ���9�޲޺�
C��;��4�ؐ�Ljz{�sXV�� �q���Op��ҭ��5&�m.0QNY+�������3!e�̸P��y���v�?��"���Ȥ��y�P+����P`���+���!���^�IЈ��i�Fpo0ȳg�Sϛ7>.-�Z&W�����V�����3�����
U��_��sNX�ٿV:�Z��C��:H$8�b}C���7���{���1wÓ˭��;�A#HKXT�+�\G W���I�+���~6�q}�=�4�S��>���@��vI�9NS���r��6NP�^%ܖG+
O�4��+F���R2��y,N��	��i��M��]ޖ�V�y�vhp��vݿ?��ظj�N�ٍ���9A�K�y��Iv ��_��:XB�lr���b�8�8�;�FqZ/�[�C"� �i�~+'$��R�S�3�d�Q2�+O�T�t嬀@vg}x}vLl�o��ٍ�V{�ޮ��CȺu�67ݰ"|����0#�!����|�҆�
�hek�g_	��}�?z$���� 9=�Y�aʴ�Z��Y�	� .�+QVR�M��+�oGr'��>p��`E6APr�-T��]��h~c+��c��l,����VTg~�y:�8(�%�Pnگe��E�NOn�=���]Dh�xW�I{����\d�.�	��f�:���V�R��zƋ>r�7�i9e���Bp!lOk���&�,/�J�h@m��@�S3���h<��a ��I�}"V[\�I�p�!7�r嵊��|
��1p2����\V$lpr�2���M���G�����s���B\~�?iOݸ8���H1���"�Y��Z�g�����f�mH��Ch#������
Ҫ��:�7�Y���[ʸ'p��B1Q��;d�?R��Hl�9!=�+cI\+�Qގ�}�,��nq�4�G�R�4��E����a�/�ނg �3��s�>UMN���騺���ZM���1^`�f~p�n�	i��=��x�[>�)B=[�)�8�:��v���H=;������y�
��dbR�$���Yc��!�,���s��Bsr&p�D>�H����	�,���y��pko^��g����u�^�M �$�\�<��m�)W_R��, ���0m�j��c�U��k�q,P`!J�O�_��0U�����;x�\8�N���ɛ�����S��1Y��12Y`��͏�^W��k��R��Kw�퓑��v���0��T�\�}U���6�y����>��m��S��A=P����,t��O��pҴ���t�I)�� `��܋)5_�P��(��m�u��?s��[�%���.U�p5�'�����z	�^�G����x]�OǞQ�>�]6b��^=qG�=� ?��U(&'���vk�͚���~�k觰vs�����IS�=^��o��Yq�H����n1�,�Z�*��4P��+����`�KmQ
C%���)��/��W��UƢ��Kd���Y1XI �F�DD���w�3֓���u��\���9/ﵵ
5nP�|���l��,iP�Z��ݷ`����ԏ*�����ff��	v�Q ��mh�IjC��o�L��0�Ou��GB55�߸Sp�ȕ ͘ C/�!,���0�v!�]��M0�~������N�j�JlD����R/2{b�}����䰹��(Fa)�1�􎜲@%"�߅r\�8��k����[Z�{?&1n�Dp�����VO�+hQ1	�FQ�]	S4(���M��O��7�M� ���9��D<�#M`@ ���z�5��Q�I��|[X�O��z2��@�� ɉƠ�"�Bv�[Ɵ������8�KǄ����^A��B���[G��W�`���i�S���m��f��kC��$?x��h!��9�x��W`��)�w�eMY�=�㡥�
:{�G�)eU�'��c��S��O�(΋�y,� � gꗕ�BG�����/A��VU��P��(�ui[pC���oLf��1�=��"D{='K�~Ahΐ;h�W}���L|������<u��	k'O�Dm�$���(�b�
^��J|�I	��=��^��&apv��n���^GlN��
�F��E��dkB 7�G0J������*FO��ޠ�(Y�^�	��:9����g����f�������$*��!�ҕ%}�?ꞪȪ����!o%���B�/�L�5A\������D��S�Z������xD�=�*$dΒ��;�}7:d�9�Q[w�tX�㥬 �͂�]������n�+�)(���k�����������5"�%��.HZ�ӑG	���S@?�c��\����Qdyyj���c<�Z���F���vP��N�P1Ϸ�����x�H�����a�k���y1�@�h'y�1
[,��[�}U��/�Ks��}��fJ��~�Y�A�;�hm9�9i`��ى��XN�R>	��o��Sz��7��u�r��cӵ�<a�n� BM��!�f�cj��O��y��崑\�=p����|�C0���2z���Kɇfb!�z1��U�D8���5&�<��������#���-�獷������F�σ��MUslt�+]]���rw�mT��]���%�x�,�1�~��c��G�1���~��� �G~�@�RR�?�n��FVj���)--�Q�B��"���[��\���M��n4^�e��\�;�H^]d�����~��c�W$#J[@B�q�b]�����$�Ka������(��B���%���Jv� �?�ؒ�Z��uWlZjU�����cA�������(g�N<��P2��=���������h:�y�]�nƭ���������g��U���z�+8�Y߀p��I���r��?�x]��\�vMPA�{S�'��.���Db8q���؉�j�Y���k��$�`JqU�MC"U+���8�����5�r�����vx�┸õ�q�p�Thv�W�ks \�����w�$��Ok����٫���9�(k��^�
���dz~E��@x �f�9d�Y$�%���?�I�_��D)�`��Z0�e�8#p�>�F1F�Y��`x8�Xĝ���z#"���2O����Y�[=�*��/�����P�����;<��Ut6�V�[�>}�X/6��[�����
���O�3vjdYф���-�cW_�"C"��i�As�-t��!H���Y�^S~}5�,,ۢ���Es���(�xn��r�r_/F��KZ�����5ٶ�,�EՈ��g~sj�hw闒���/���'�v�>�mw���xyY�X�e�ƍ�`��B��ڬ�i���c'߲���^�K	��)�V�>QR �55����H���l�Q)i��,$ɺCl�� ����^�럵m �`����$,���)��P�R�����Ƌם�00&YR�h.�]bE3���K�`���'�UKg^f�}�T��ܮW�g֨D�<�Гq\u�X�]�Y��V�:�-�J�b��1�3t3�kB���o5�
�˶�(�2�YP���<��X�	DRU��$�]� ��5g=�J$NI`ZǶ=�kva�7��;�nQ����S�X��8)���b�s��	h�=*e]Xg�O��1@�f�0�Y-��������:G�C�kZ�7箝�;�)��k�J ��ǳn
m 9�^�Z{�!�|m�'�ۥ�N�ݺ{�����'�T���qXB�ʖ&�D:~���;��ln����-�a��lߝ��uq(��;_�E���|�;E������~�6�wX�5n�]U ꏅ��8��+Ɋ?��	��O"Z2kd2P-���U��m�#�9)�����P�[KUq��ҿ=~�:W!>�X�*ضJ��9ͫQ̬�s/0Qni��7,8���1�q�>V��U��0��(Vpa6V6�Cn� ���I�(XC�����P���K��S�b3�^�����`�,������X��S�i��uLK��=ƺ�W����$?_�fB����� }T���v����L%»D�&*FYW�0�(^O�ۢM��i�_��o��!��6��Y�\���z4�Ġ��T@K�0sI��H<�\�s-��އ�� ��(�{/~��:����M�Z�*mw��P�5����0�cYח��΄!�ɛW> �fsh��N�)lA]]!
l�dm ��}��`�_��
H
~�F[�`�J�D�||�&��_��dH���j8C��D��A�Β��mB�8Z5�u�tL�D���r.^R?x���������`B-{o	j���R�N��|�����ݞ�n���4�;O�jͮ&��pV�`
��3 lWXl�A[H�����,���A_f�:���+)�a���� E��A�a�-/[�>I�c҉��wq�s�ͅ��&�<�L���Jx"@��6ȟ�{F�W��� �?%ltH%���`1�1���]	A����'�Cx�t�Z�~l���R��@DF����C�ń�p�BM���/���-��������21P^�!�F���T�����!�o�ĵ�»:�
�:B"
������c�7|M�w����MuDd�NA}��Hst�����Y�D��[LN׉F�΃��?X@�)�����1�a��Z�XD�/���͢Q-8���xG-�����e�t%�����򠸭�q�l�vO��t�RP�a}�:��2�"�7xQ��n鴗���!%�8�wA���l��ڙg�/�����y/~˟$K㍛�Y��.7m�	.��*k��GC!�����R�� �h��݊��2�qI�:���nd���h��x��9�V�^	yg�䔆��ͱm~���T��g���_��J�S��8$M��<�N¡�3#� ݊���hհ�P��Z�:���_�E�o�&%yʤ�Nl.X+ke3�ڳ^	b��.q�s���v�����t"?ZBm�n��2����¡��}���́�����v3�zsmz���.V1�}#Z(�+���u�8��#�} �xX�e��M0�1>�{Ƹ�h��{<�W�JZ�D8��Q��u:�90e���Q��xomo$r�ӭ�~����{|����N���wƝ�y"aiz���P�h��.Q3�2��g* ��c@�$g.�$�<Jy|M�F둖�2�!l�#R���bL	B{"C��{+�HR�8������;���E	}���O��t�]�H��B�|��M��΅e�:�0�EvD��/����͚H1B��0��lE3
$ԗ�@�g�a�����\��0?z�Ɩa��v�oo���D4fH۝�)�=�>��7dI�׭xRٿ��<8��,g��u�)m;W��Z��!;����	hIgס�����_��e�ix���_
N}��J7��qa�����l]z��p?�3U���8��^���ظ,�x�s�d�
��>�3W��p��2ߦ��R=�c�7=b[�x[;����[E���lbCt=o�/��D�� ��j_m!9�8����v��!���Ǒ��-���u��OW��j��d��𸜨:�B٪�,�����:��+t�Ӛ$#j�j�岮h��#���Y�T�E����)�8IQ��Q����4b�W�H	�r~-��2c��8h1�mY���?�5xq�;�����.^EO�i�r�f�q�XT�)i!��x�ƌ
�S#�5�r��d�6�'=, s,��V���W�U�D�е<j�����L��C�a@�]H����&Eki~q��2��6W�o Z3kx5Խ���X�����cXg*�K'��������/ws6����~i׵5�*����C�R��Em�1��i�,����"�tu���6 �x�.�t�P��&
�eb�l���N��N���Y�\�Qf3I5i���$������L�Of�q����`�甦v����9��!�W;jn��$�2f<���vf?a�W��rră�c`�l!:��{��L+��Ql�R.��]��K+fR5Ն카#����������le�m3��5%�e�/�>�p�ؠm�R��N��u���`��l]��Jq�	�
��ʻ�s��M0�v�ίFS��a>/o����D�m�G��Y�fw<��p�B͈�.��oإ̊��)2�7���I2�ZN��'+��2��CVxU�g!�ڈ�>�c������B��@���C��Y���3��p��fڝ�Z2zW`��>����ը�F-Hf)IAk&�`7I��b��E�8��Hlor_�� �����ܪ��~�κ�JS��ݚ��ϒ�q��U�J���!̼����`<��W���Yr9�߬҆�v��Cp�霗Ɍ��82\'��o-�m=�{+P�R��5�� w��O�H��*IJE�rf"�vU�ԋ8��qZ܉2�E�V77o�iN�[ܩ2"lab��Tv\B��H+3g��q5�]	�(�m6���R�K,sT�0����؋|A��^�6Y���z��?X��=˗��"A(�*��E%b��:��x÷���M�F�N8�U>�i�xw�H=l��$���ѱa˧�Ŕ-�ع&s7�!7'U̥�Z9��g����~���!X��ez������I���7FZ��*�����[�cB��@������s���dv5�V�i��@if5Z���b�����Zr"e:�wӈ* "KZC����M��2	��Y�H@��E�6��ō6ͭ�����b�Vg�"eT�3@�.�.o)e���Ԡ_/+������a\N�JG�
�<j��ʴ��S��x�?3��ޕ7�(��x�G^t ��L\��p��vP�������X�4�!�ا��G�#_02�ϕ%��Y��)�/'Wi
&�W�Bэ��5E޴�f��{̈�#�wtٓ?6g������8y_Ot5q��bE�<�I�d��|s�/�7��ұ$O���O������Q��(��t��� }'��J�٧�˗�!�Bdz��&�5�*x8O�s>[8檷��!x�d�0~R/�w�hrZ�d�y��B٦����N�[yaa�@��^R���)�L�S�����׼vbJ�)hA�ˍ�J�H; ��p�~[�
��	��x颀�6T�L�GM��X)��m�>��īMӟ�Z�KV��f>��r��+��J�ٓg]���i��u��\�����'�pC��^����OhS��Z�DC�k��`2�]�w�_ǎd�.�d]4.#�֨ۯ�2��wÏ�D���[%2耼A��,)ȯޗ�#���79R��w����ڐ��z#-�\ћq�����"���C:�w�^,����j�}�~���-n�?T��ɶ9�5f�g�s�X`aIb`�a�I
\�9���⓯��D%���Z:a:W�wB�H
�r�12��'�cג��2n=�)Q|�\}�j�ɕ�~�����`�g��#�I"o1���q�4HP���;3��^��ϱAOA�C���Ƹ�'L!7��Z�."MP���5�����MVde~t��ە�C�2��ќz�Z
f��#��QŸ�![���R�C��ـjA!���]������KH��H�`{��*R��w��_��B�t�Tke�[|�>n+KW1��xXz�@��Q
:����d��	,C$�bQFz�N$_L�EEBp�����n��.��i��(<���K�m�͊ޑiÌ�;���7�~��s�z'��[�wO��Uc� �.i&��Ε�g}�����]�ݚ�VlF+X�ݬ4�U��]�Ox#m��&q� 6�R�rUO~���.�HY;��$)�q<��-Xo�<�pab�'v�.����`ӗ*��t[���p�����mC�j�J��_4�p�r5\��7��n�/d~��ߚl���z��=sݙu�\���|מ��Z�q��ǐ����X�?4�T�g��ݷ�N�[��+>'�@�n�n�TE�z9�T�-�PO��e�3%#Q_
w"�E04�qX�ȋ2���KPu�����U�� ��J��Ym�&?���{�i'U	��ڗ�3����d%��t6P	��i�xج#�q�$�ο�Z�4L_�|�dwt�X�g��?���B�jD!��n*_I$2	�jM��C-�^��f�PW��X�ٓ�!�j1r��kv�e�}��}e+H<� ]�>����Ωy�O�^jO�L&�1q*��}�v���BB���^l�׋ƻ�gջ�t�rd!�X�(��<���l鉬[��{��	Kg�Q�4c痺�3A|�6:��,�-,Y��Dݐ&�^WA��&��^zr�l�1���Ke~��|j�ѵh��I|ɱ�o���X�tu�7u�Mcb���aM��g���F_k��f�C̷���,�Ռ2�hY�)��!sM�0[O�1Rb�m�"��S�-�1���,�adT�p�̢{`�4�����}=K+,@��-�u"X-��nz��6"k�*�v � x�R���n�p`��$�+���U"��=�P//?�{\�P�&W��*paLMP��C�_uc,IB��n+%�2!*�$�P�h�G��QL#���[��u��X;F-�o�7����QMUU��TaKG,�wLÊ���D���J���#�fb�M�0.�]�7�^ �29B�.���YƸ��8�]���ނ���x�a�$����d'Ћ�W'�N�=bF�W�S�@�ٟf	=u-"��S=vEՏ���|4U�5$�2WYЖ�3G�i��n�<���2aDʻ��3�4���v���}�:N"o�N��(�nު��� ����m��ڕ6>L��l�M+�̟)�J"�W����nR��f�:��<�[���[>�9Q4O���c�6Y3�>��Y��U�2�G�U�+�U1�_m��tv��[��!<Ϸ#��-,�����$���ȎPـ%���&"�7�I����	�*4�{�V��{����3�Ի�0��3�D}��hM��I�B���w���*�[���N����g׳!�fia$��l�x��&&ڶS^O��X6��Z�+�׭
���+>u�,Ȏ��(���F����)�x��K
M��멐:�r�0P�O��������;���婽�O��udm��czr�<%Q:�nicG�@^��>YX9�Rg*��O��4�i�D�:�\G�_�]��U�D�8LN��ڜ'���j֛u�j�� �	Si��� ��`�G�
ŞO7SՕw~�Xs���#�uDOA�����Z�\�:śS��V`��Ļ)NO��K-؀B�;�*�Δ6lXr�I��ﯙ�i!�j9Q�#QFwlS��e��	�1FR��ݓ�_x���B�,3��i:�zϞ�T�Pe���~�A3�C��T�'Jb�6�5j �L�ưI�ojn��������${c{d���_5��KT�'�C�.�9��q����iR3�]��F��W��#��ו���m�S�f�[Hv�jV�'5֌��?g��Hh�/P�Ⱦ�yo�<�`:�h�BJ��,M�qW��q��|,��sy��-���F��P�wn#0���5Z����&�$���[q�]�h�dBCP��"�C8��I�o�Y�f�Tz�:(O8M�1e�����������F<
��jX�!�^�d�u��2��K[m��luL@���>��~D���PE�����A�gJ���;*��,���ߺw��OQ�X(�$�c��0UۣZ9T����H�n!Jts���f`>�2N���v�<`�A�7� �(��:vk��5��䭶K�L�r�Ans�N��X=$��E�!X�b���R�"������!a�p]��ԓA�a��>��Ñe%���Z� ��A�p�W�Ԏ����YS�@jc��M�Wf�L	��ӢV���V���[z�17�d[�%z5���8;��a��^�b�W���Db¤�1с�оƄCG�!�e�u��
%�7#�.*�C�!�=�o�X�C��6L�PJ5�ߋ��� V�.��y�L�+e`l�\��w��z�6h-��*s2�,��شu�vh�8��[�&"�r%�� ����d~�-)F��d@Vs�ܣ&$��Y,Ͽ���Aɽ����Em�8F��b1���d{=!I%���F_y�̔�4<��H�����i�XH�3�1�J���l|��!tm$Y�&��X��T��>���I�L��}g0�E�|��i�=��Rȱ���eh6�����j�[P�n8�����B'�U4�!~�x��6�3S����^�a��˺'i�]<q��2n|;V�WD~��b`5]��ա=[vU���-�t=���V�qC`�K��:�*�� 8?&�j-[��s"�1O��)[0PGV��hY�!(�X�]�	K�s���/.p�Ee��ӑј���΄�ԩ$F.��Q��0UU3��Yw�C�D)OeF�g�k�J>z��ȸ/L��7�}NgRS�����}�P��%����5E=��c����m�i͠j-���/����y)�����9��
�q]AX�q�s �z���d)�{�Y�W0(���P�-]N����;v?h�Y��`���O�pn�jk�Y9���|/�p#�-��Qxn�6E�J.�䦱� P���P�HqQ�N����'�ka�N6I`.(�˛�{ʯ�.B�|�m�bV6��(��
3���|.11�������O��#5�߱P�Ckm��uzv�h� �T�o2�$�5@!z@�;�?�\=�N�A��(	���!��ֺ��	�$��BrK)9����/���aD�B�B���B�#�#
�Y�`�f��^�{��t��K���Y�b��c�z&�R�Y��xf9e��r�D�M�J�((�TtmN	�2�|������Z�#���)U�h����bS���]F��8}/������6�7������ɍ��?7�SFς�h/��ږT�A�̪�&Ɖ���B��=+̭}3�[}s�1xY�WX"�(�#�j�M>/��&qI@ݷD��8�A-Q�<���T?:p*ˬ9�?�	�ާE���.H���g���!�y*���a`��X��&;ZT7+8�N���3��K8F 7*I�C�t��^9ui ��;�"Z��w�^�V��X�Q���!��O�p&�E���P�rzMc���p����]ќ+�<|�Iݞ�R��Sn���ݻ���b��Sp�_{�ߪT�z;��
mИ�,��I��%�\HM��R,�@Xx��J��!H<���PUS���(k T���m`��dc:��	�6�9�@B�7y�y��]#�
��,b;Q��j�9zn�� >��%im�p/�'D���y�Ӓ�HD��4Yt��R���+1��?W�y���w=�"�B7��۷�;�H��rMe��#�-����V�Ŭfo�⚣�w��������򤟹;�g�EFDaH�[� ��=]�Q��Bh.�� ���j�X��p�@r�M?�,�Ľn�������h#H�@c��rbn���*_g��;�WᏃ:0�Ƕ/HشZ��2��=�,h�0�ۢ���%�i�	�y�7r�/m����p�1r9��2)��7��v���n �4L3I�䍳6 ��ճW��^|An��`6fC���w�E���]}�6ݞ��jk M��I���������Jg�
�Bx>���������0����Q3H�dtؼ�K����6T��O�WEk�/'��F�ͪ M@�0���N�aA���;�T�ma�Mv1��\%�����WWb�At�.�/�AJ�z+W4Q�[LK{>ܐF�c�̲W!Aj�̇��Trw��U��"�p6��@�B��HyFJ�ukGZ���>�-#�A��P�fN���5Pe�-���;�_e~�ն��c5��+m(���t4��X���o����PPO�$�i�I�:)���o����*7�~��ކ��P��q��Bߜ5�Z��k@�0g5m �_��ݔ/d��cPE%���×���|6�/ q.o5���jh�HY�FJ�_��b�72��S,�
K��m-wh1#X�8�V늚 T�o[���pK~#Zy���f܀��|"r8��<в�n������g��\����J�5IR�x�!�d#��6�̋�A2f�FE��S��;2`���+L �!�����U�VV��vŗxV����%�v<����z���N�#rOK`�+:���orG�D��H��Ƅ .���N.����G鶘��"�؇g�FP��B}�����Ӻ1�h��������^7r��XS�Ԋq��bv����A˝l@6K!�on���ۥ��uBx�	��-�/j���x�S�bX���J&����@����;�~ri�~����a\WЕu��+c�g�mʏ<ᮊQCqN�)��!ƾ���:� ��'!�hJ�;�ִ[�@ђ�D�?m[+p����B���k 1y��lq���u:=ZjKJ�_k،�Z����/a�[��?|���jKT�Г��oƫ�y��z�G��]�
�uu߻��ӥQ���C)�����*�3���G����йИ��r�4�r���ƻVJQ���̇�r�za��	�e @ǻV�mX���������Ӥ��w����Og�ή`2�Ukd�����K�L�C��C�[ӑ���U<$+|��7P�I<0�0���Ρ@�q�>�2����Ur���ۘƮtǭ�������>�{ak&_����[@�
�g�m���O�"�U�6A�8�W�
�j�G�r�iG�4D���UTp&�!l�GfAo6��nO��{��Z�o?����7kĘ� Vjo�>-�/t�!t�}�}��!��u��{�o_�A��w�;������ ��d�Ƅ%�E��<�i� ���=�Oo 1���&�9���e-��f&K�iw�ង��`5���f���՚�(į����1[�n�{�^�pb�E����{�K����Pi�Odì�(&�D ��71 ��&���ם���.J�2�)���[~9����)"���Zx@s)I�to��9x�m?gwc�������#����4T��d��)����L�|�Ϸ�2���2���L��������	������5IBo���"��z<�C�"��,�����K�၉�UN�UҀ��&0ɾ��������X�����c�Hٗ�$c�,H"�A����KP���m�xd��ľP�&t*���`qYW�)H�Ȁazᰐ@z�����V�%j��p���a��s2�4��;}j���9y��B։!�DՍ���ϹdݐgX%��tT�����$2�:�+�I�)Xl⋎������a���pɡYp#f�`5>�v�ϭ�H��u��ܜ��|�B׀ؖiA�Nwx~�,d��U�3g^exz��-{q\�F�j?�T�s�I4L��F���:���L1ߖ��U5\i�X�`�����5S��x��A���
^��Y��~���X���)f#]U�׋B<8���Y|���-ci  ��]�7驫��抪e�2�����f��D���Ϟ���r[`P}f���z�����+�w��y �!�
Y^2�(��k
U�]P��<aF�Ue��)g;���*��2c(���r���tK������?�ɱ���xw4zճ(T����,�p}�ū#x���և�����q�����Z�K�4"6v]�x�0�D��Cp���@r|�I�֦�8����GEo~(���v����R�FJu?��G�^[��P)��<xw�u� EM�Z!�糷aK�D$�C��epl;�;w4���j���\,�*r� �����mj�qT���Z�"����+�ƫV6�b�K���4A��z��*���_`ޜ��X��X���9욼:����Z����=��Q����30�%������D�wH�:`���p=B�%,#������������ C]�Qo��X��e��Ė)h�������lC����RQ���C
��.A�WYgF�[)73�J{�c��"��q��JB�k3{�\	�eo�Ÿ�%����,}���������%�ucu����Lo/�����}E�����T�v��F;����|��o�\�L��;'���n-���R�pxh>���s<iP��$�B�n� RkkS\���浧��H2˻0�-��(���`LEт��X��mw,���.�[�߲���7�K����~{v-7bFũt�󃀐H�Z�?�<u���=`G���&&\�-�E�ua���u�UC�����{�h��,���h�.���[��xw�%�`L�4���_�S�_���2����)�����U���>uv�����+J����y���r�5�n�j��BI�ȌS�Y���<4!V�'{{����gj�h:���)�Ro�����ˑ������<!k�4�Ō%��N��`�XЀ�;�̜��P�-�B;@�bυ'bն� }��lz�X1���k�/�U��\wp�:z���l�l� -���4��K+��Z���'f�c&�
�ɹ�Ƒx���t 
��U_�Uz��q�3��^���\�k�hejt�s���8����E�`F�;,����PL�;�n�H*/��2`4o��֙]?�y���>
D������!s����-B�MK\�%���;nW����"���Aۘ�,�_���aZ4�!k�G�G������]؟�$�D|����3)�.k��_�W��a�b�N�
' 
��5�)Ȼ�p$��`�0��_�+��#��YG�X��Ú7�	�� vڲ�=>�9�ב�]*��D<�`q���%瓗i�a,Qe������n-/�Kc��r0�v�E-Bʅ���Dբ?'�Z��ab� !��A.�U�c5�u?3A�؅h�6Q�Ỷn�u�1��d��6�0v��[97-�L���ʹs�`v���i�X�sy?��K捼2F+~�Ƅ%��b'���#C=_�Z�X����p�Q���z)���dPǎ�I���=>�p�Q�n�f\�.��I#^���CeL��h��q�$��%��CP_V~�Jh�]�@�xeإ�{O�},�b�L�:����MZZ@C�K���΂D�2̸�����[� tk+�I�k�Թd���;+��ˑ��7�cs��9!��IѸ9�M/�'N�,�	�˱�����~r�H��H=��t�n��{�>�љiV���KySA�7<G�����П��A�Ž;A�_,���7Yt�B����7`���ͧ���Tp!�<v��hn�l��\��b,d|�R���wH��N�p�b��fby�p@����4����r畷�7�I(-n���y��*~�)�����w"���=� �����-��RGt��߆�j@�mhtX.�#�%Kp�P�� ���[��8/��Z��ْ�$L��ܤ�'�c��#���T8Ob�..E�>��E�	�\t�'�\�mz�k;�;�{�#��+b����|r?�y�E��_�z��0�ɨ<bĒ��ox���qY�����^>{}$&p÷�cV��s���i��ڟs:�ؙI:�L#��	���L�|���^�d�$5���:������P�jV��1Z�z ��Ch�2�,4x���^ʴ&�>��+��7~ ��QK�Z�ޚ����;!l��g\�x�6�ɡX!��X�Vg��c�%�BU����yqw�qF\��W߱�޼���� �S�<r}4Jݺv���d�07_��-�&�gO�чTޣ*�n"\¾4�Z��a�~8,���W�q�rA/7P�SZ��k�m�N^/n0F�������������2�2�0���5Z�Z��+�uj;�������������_;0�����OW\�"�M��e��܈�t��n�)���뿖�i0U�Cٷ�l/��!s��wN�~�,d&XՈ8�_�2�z�,���4'�!��j~�
h<X'���j�n�FH�:躭�p����J�F	D���ӧLB�
@�8m�2+��Ky&y���=8Z�A��!o+M�6$UF�iB]p�}>��(9�Xy����DԞsL�h��b,������c|��v���:�}�v��c� c�o-�C5�ۀ�������;O�2<�W#R!�����|ّl�w>D'q6k���I�E�tr-Vu�����}j�\�-e��j���1����T���V���#�P}�Z�x��S&b�`�2�P1C�<d�E�(ǋ�-ݞ����crd��;�e}$��5���	W�{8�aZو�𔈩M ��BE?[��}���!���\W^ Ek1��,�;T���:���k��:�"М��K�e����� �1e���KՓb�Xl�#~�X�}N�Ѐdu�F���q*��;�Nx2�N���~|��EA���^��N��������&�j<�3uD}�G��6�*���$��
�0�S�j�nX�b{�Gg_��t�<���ǰ}"�V��G�x�>~�*7ͿsD^j7�]��k~F=:w�!�^{�@���qg�������Zg�=k�-���f��Σm�ro�y�g�~����[�5rN�ϥ�qIO3���b����-(��5!�c_L�Tc�o��k�P�a�f>���~�o.#��a��Y+�*Gi����н�#\�5��C�c��'`)n�O��Pi�%�qzﯤr�O�=�V��n�0�x���Ƥh�ha��&y	����?/�iܲ8��q�^pM���M#@����2h���A�@�{�@���:r�@���]��kB����W7�F�1�@���{Z�Ȏ�קR���%4��w�7��+���M߶� �%�9%';��rĂz;�Qlj!*�W��oփD&By�S������������q�j��f��i�p������`�����w˸c����9HD����aP(��w�5��C2��_ynC��9:�{�z�Y�E�F����j�K�2��QWm�L� ������)�'oE6����ׅ��߁��8�2ݬv��
����q�~e�9����Z�e�Bu��$ n�0$�ؾ}T9/ŻB�iMI^��a��v��n����oC),�k1�" ��O����C��mT��t]�� /���@�g��z0�U�5�A���ʖq�v�����`!�|J׾'@#g��fdr��NE:𰚗�WKs��<,r�x�� 9��c�:l�A��(�f�A���dT�s϶�:ču:{���t��t�G�T�4R�?�r<���?�U���[6AL�٘k?�]��r{���'�O���O��0"�:��e�Dk�9�N��!�j�,���f[yZ��~��[��ϻUG���9�΄5H���ݵ  
���vj��j�?M�!�q�t�]�D򋗍�}4�'��9���L�m �=��r��[aA�Yt��C`��<g��t�/��2��M��ta�s��?���-�'��v���̈r~a��	�ᕓ�Lx]��,25�oe��A�uY8%�RǛq ��G��Fh���uO�ID��r�ߟY��~�?7rU��JU��kU;T`㝾�}O�{��eק���=��n߅��
��74�KB_���Z�K��~mD�JkDÅss5�����(��%��Z`���2�(;��S��t��n�����AؽZ�ճ��WŃ'�ȥ�N���y6Aԛ��yˉ��Swe��o����C��R�V��E���l; �u7��lzK��+ �1�B��dJ=uO�����Nq)���%�P��_���"�.�Qt��>Y��@��Y����z�$cԾ�b��sV!�u��&u��i�J�v$��U��J��._��I	�
Ӫ�LQYbJB���o+�(��=� ���(��Dq���p����175UcR�@�Q��W����V;��	T0m�+ ���EBh�RJn-\��{�.X�Eu�6���{��[H22Ȉ�F�JA���v�;v們-����T������dj�wT�6G���F����uU�I�'��v��K�}�+���O��{V��Ŕ�����7��%�ݟ4���3hz�l)Lū��&x���!g�t�Sj<���+6GW6�t��\��k쫰�Ua���ON�ݳd��$��ԙQ�c
9�31m!q�g2S/�Bŕ�� ��0��r�t *�	��eB��Σ���W?}��˭�+^������כbS|!�@]p��ux�%�/�L��@$Bz6w��r�f�?��oїLH��d��Y#��7���ޞM�*m�|���YMhm����S��hn�dՑ��fL����rp��y���ߤ��U؃�t��F��Y���F�G��P�+fH=|�K�A5�i�u$�ګ�_0ÿ���R:5�#{z����/�_~i�#��)�8�L�M$_u�4���p�E+�o8�O+�H�!.W�B}�z`D�|�il�wL�
�%����F���Ҕ��K�s{'���v�MA�k��5_b����'p�yyrc'_����3l���$�?�����CgV<&�ד�X�VD���E�u��8����#��q���j�k0�}[�/@��rgBL�lm~P�%�=d����0[jHw�� r�*#G�f�#��M��~�3�A�p_���q�5��k(�J?.�w���U�INV���{�L����ZDG�W�C�R`�{���$����b��D<�-�Ģ��E=OX���Ga|�#a��l����GF���"�ײ��C]�#i�ӥյ.h�]|�c�g���U����r�ξns�D���JbP�GL�?I����@��`{(^U��䩴R}�&j�p��!��\��N�J�0��#SN�Q�99wW���J'W�����}|��`k=���%֒��nsD�c y"�1�%@�B�&�x�����0�˚H��T���S�gq"<d�mo�p�$��/l�싲�5�Td۹QVBȲ
��:��%f�\�ܠ�!���쟻|���t��{��O𚺴�=!'P��h,��Ǎ�ݕ0?�9Z���4+�ǈ��ʶJ���gk�:�񰱿�FKwu�/ZK��L4>r�{�"J^����Ǖ�p��3�mz����S<�+���zWPCA�-�q��I�d���0o[l7����6�vC6����-mBz{f�6�&r�&2U���8Ϯ����B�`%2Q���)�_��A7�YQ0����&0裈8à��`����;խ`%vf�Vɻ(��=��op�Ťp�dKl��Ը��F;��F|9s�Q1&~���$f'�B��q~C��v�n2���J�4i�B�B�Ŝ�(�PV��F_>�Flq0��X�<�;k��ǃJrD�T`��c<��4W��9���(�[�f!��/�P�D�����&�
L�)���� �jnB���%�����[�8)��z�ܐI���˫_bv�0Q�"�r񟯂���H�[�H��#:_�D��`����j�!�Յnq��c�|nk>���jΈ{>�i˓1�w��	˱[+l�����x:M�8��� ��U�?�a�*�z�4�)��䋙�᭕�c}lC���/SB�����M�M2m ��fYօ�����3���u_�Ym��~nd��]��lȦ�e�\c�x~ó��u��x�E�V��,���T*)~b�-���za�>�	��l��#��2*<�P�#VDlHvܡՔ������aP4�1���<7S���I�!�i�qD\�P�M</o���K��"jtx�e�Q%M�V0X'�9��H��T������\�5�����?(gV\���� �����r��"� ��]Zs�a�������,Ǒ�)�q\�u�O�R����K�����v��>���ӽ����[� ;���0�ZJ�4A�gC��-v���B�M{QЊ�dc�t��p~HMy�q�/� lo���>w!J�Th�8.]�Y��+5�>��5!y��gY��	~���7'��������S_|�G�e-ަ��Ym���]:[d@��@�t^������O�RraC�t\ ������`sdOB�AM3���'�3u�/d�`ط�Y]���7�ƕ��p'_'� 8_o�/(F�c�|Q���=�G�S5�~�>����;��ZuE�z��
����$�͚%�v��\��6��o(��>�z�?�'�v���I�|E����);��U���0����;,<=�vS�&���Lw�J~���0\	�ע�^�$��e͗?��7SY��)�B��	��W$>�B����(͚�"���9�����b7����U�t��w-�/����K�O�J�T���
�u�̙#�a�;�ڐ`Z�ɰ�}�QZ���N�)2�;Sv��x�(���{����5�&2���x�bZ�M���%7���Yd?���Ȉ���V�./BLX;3�6��[=��F`nX�+�0k��������$�L�'M|�u)?��qۀ���u8���0���n��⯅s^����cp��r��x��oK7c�����S�%֚%`���V|?z��Y)w��Yx��+S�d��Z:�pj��(����"���T.��u��W��Z*E�V�O*fK��S��M���wV��z��!�W�^Ni�\�b����A)'l�QS�h�M�<��-v�غ�($%J`5�4�� �ݧ�q��@��cN%m�-^��;�������
e@YS��B|���zS������}��0:i��d(��Կlǖpf�/Ò>x��s�O������B^f�fǾr����Mya��V�ug����8B�#9p�6��u�9m5l6�����I�;) Jb8(Ra��=�$o�������]�V,�,(����b�DZ������iDl���>&��k�� ���9���O�-o{c-�+ w7M�Nサ�Tٚ렟�s���3ٺ!��9��mQ���
��쉒v_�X���~��Uh4�^e`�A�~j��g��Ԡp�M����s���5�����J�m?E�.4�U4�{�p�b��|�lj����=M�WR�/�(���ݞ�e���R	x�G��t�!sK.Iy��'W���.��o�ɗY�/��D��o؎G9b��V��"i��t���$���K0?���n��$w��ҽg1���{��6�u��$���	�ֱY�Y���8�X]<�C���w$���c@���W�D%�ɟ�>.z	��#]�{£��+JaZ�7@�]�0B��1>�uIP��k��.dm���N�פ�du�I&Tn�ˬ�1@�o��g��S���d	��rT:���7���� �OP�5��P�`�HN���f�m�/i��
����Z���<?)!!��/������7�s1E?�E��[rO�J�܎��u�$����X��>5 �O�D��GƜlEe�9n��N)p��U�G��:���k�tn�[��P_�z&u�����M���n���5X��[�C��닁��Hxw0`Ǆ���M�z(}�� ��R�l�ʻ�8�?��|�����a���No@���X���//�b$jO8l"�1�F����̱`�ߗ�<q��i���q���sZڼ�sk���l���8|��<�/"�ǚ���f�|$�b��l_��,��0��X8u�'��@t �<�-n�ihX,�"}��t�-{��p�ȵ��9��i4sč0�P\d*�>�UXTm���S��A���"Ť��W`5�d�0�g9��2,��w��*�<�Zv��tr%Kz��r{��������Qd����"Ӫq��
 �[�BU������T���ވ�aS"O��B$�G(�s��O��/�d^q!�;&���>�2�����e�������#D�~��l]2^n����W=����W>�NO����ݏ�h�d{����:�>�����3���������@��ż߀B�a0
����\��i�~P�♃VF�i���D7�[Oc�O���B(�������d�]Z�N�n�ہ�{�ŧt,��������ȥ;�|�M�|�d�������So��E�0�#��=�5U���8X�sZ%Q}zC=hE���\�!�W�㽷Fd}R+�¡]'��*Ǵ޸�H��ڑ��`8a�r	���aV>&��"�����Ql���hg3t�h@�E+컉�z���.U.l�ä��=�t�l-��� c$!�����Z9t�N��3ƽ�Q�v��rrK䞰���H�`u���->VcM/IL3G�ŊJ��r���Na�VS?�/-Bg_�4�A30���H�gT��[,l�iOQ��(�½N�=3;�C{tJ;I<��Ow��\L�a �R�K�l�P�=�$�Jad	z)d� �B���Jܷ@���/����Ae�2K3wD�ژ	N���D�&�sE���Z���Dce�hZ ڌ��TH��C_�{r,zw2��x	�c�L���y�ĊrBR��S�^�&f Z��U��~��І���`��u�r:�!�x|@i_�U�Q�HE���*�˨(�1���mpI�v\��Z6�I�ʬ�fWiG�q��h�Q>S�P��:aV֮���)��s!X $}�O�)MaBʅɡ������-4�&��V�Dl�ؗ��Y��0Ƴm���~e���u,�,"��v���e���M+,Q!RM��%ΩbrO��13���p�[�/Ux��2g����P/Y:Z��(�}`I�}�5zxL�����	�޹�a�X��-��9�����Q�]&�+� �����"�8+�C�Ԝ慆Y��D7�:���7Ҝʩ��f)�4�S�"V�!��&��X&n����hx�u�L>��=�$��y�7VDS	T�	���z���ĸ�Þ�I_a�uT�Y;�j�Y*�D�2�Lo��v?�H ��a��~�����
B��D� �/���9���Yk�Z�Sl��L�v�����\.�x-��#��������,x�@�}td���k������s6��R���G�@�0�DwM��){�2��W[O�V�SD.����E��ҟ�����̀�W��nh�W+K�������RuL���9J��%���?��*�y�4��Uts'i����2��z� #�&Fޅ�rC�*yh�˖��
L/�/33���&���S�:��/�1�$χ �Q��?4:�s�Ng\.R�`�-�9�,J�o�S�G�]�֪�2P>-;̬~�y%�Θ��h��z��{�0=��i��_�+��ӲB�kW�28���v���,��e�7瞁V�a	�Vd�V@Ws�`葁��,Y܈Ҹ��l'X4�bv�7_����+	rX�n��D
(��C�i�1����Jɦ�P��_(�P�AS�-9�3�j�ȩԵ���e��E.�gv�k�7j�oF]@�	���ɧa��oT/ys>U������5)u��|��Q6
�V|�%X������A�(��X��f��:�Y9G��:C�X��B
�8�{���#��p���4}t�B����:ak���\R���&���I��c-�,�D�,X��z��K�[jTTL����f�Z0a�洬�:��e�ɠ�����f�*��~�H�|�憇�;AKX*4��Hz�q�B�ܳ�6'>4�b�����z����eh��
� ��4���1�®�ͥ��7�7(h�4 ��-�����_Ľ�[�0�$�r`�����=а��RV��/៩i�6�Ә�KI1�!}�}��N�%������jw'��Jg�\����5�K P��_X f��Ol෿-
)���栻�F"��O
yy���n �5O;��<n�������I(4Q���SIښ�&��"���cͪ�_�ϗ3�9카c�=�^��+iA�����A'|�3�*d�B,n�e�n��/��yX�dՂ9!e�u�u��Fc��W���0i3���Hy~8柺���ڝ�3��� u��=����*�`}|E��h'����K�l/��[юh^yd;8�A�+�:����G锢�^9�"���κM	l̽E����8g.�����~��[��y*��3
�<�P����I�hI��A��ϵ3�����#�I@�!;�+�O]�g�-�j/�@W�R�;��1���q{���y�� ���US ����ў�Lk��͑���b<�;�S�^%q"������A�N�K[O�W$�a����X�.Q������64jCx�Q����ͩ��,ǒ�D ����v��s�n|^*���}���7�T�󂤘F^-�8� ��.(M�QX�dIfݡ�z��gTL�^_���G1�?�8�t���4�����@�I�=�nuE�)�Tz{7�F���Rǜ�mhD��l��8I�4H�K:[|lo.���RE�v����?�!���������q�^X�{�v��.2��yt�xP۠���A~~x�H;s���9@���C.�c�J��3p�,k�QCd\��eS��$|�c�M1�уv�z�nL�'�h�����qջ\��D��w�GE���t�!��qrn�IL[i�Xd��q��X/��G`m����߮��:�Q��d	�jU�Εᙵ�����mM_y�6y��t����!
q��:}��y	�LF�5�������]suN��A��V9J̝9�+�������Jg6'����#�)�z.k��|vQd�:ד6Fm|����1�������ws��V�]=��.�	�k�ٮfÔƔ�����D���%�g �ڥ� qs�[P&T��#��TL����K�A�Yz:3b��ɟ]�W���Y�	�zJ+�Z>޼T��N�d8r�"��.O����{�a�Pa3"�m`UX����a~�b��6����0��wK��CC߄v̶�_��v������(��R����a	�x"k�� ܱ@��A[������㯔oA�:]F�@�*�^�z�(Vyge<V[.�&���� �=�R��q$�C�����u^���k�Z��sOp$�]ق)u{�xQ�L	���W_l3�iޓ���/�;�|5:�W��\�q�*v��ב>r�ò˕�$ٺv�6u�s���씁�m��f���1�t2�D�K��o�)����S4:\�(�_o����ە��pL�b��џd5_�|�4<��HpE�a�Z�h��t!=��^dݟ�Z�r��`ɾ`ť��-Q�1��ϻk��i0R��P�l|^YS�������a�	y�����q
6ҭ �ϰU2B1pn@l�`�(?�=�0qZ����q��S��*!N%���� P�IC\���癖B�84/٣��Ac���p�G}���$D�9՘Yj�x��Yg(�~v�ײ�ՄdV� k�:��M2-k+1Wzˡ�B���ͨ�����ɎI��1�~9։ߪ�h����ސv\�r�.$$1uc} �����ǔ��d�}�����@U�-�8	m�g\�4]4��mߒ)N��,<s��h��* ����`��矧���r��"J�
a=u�K��ؿ��;��gQy�^�m�l����^V�M�Rٶ�<�ֺ�{"�79�	ob��}JE�x&���=~pg�(~2�>k���+̩jp��B��w���T��Q�S��
1���w�3`�P
�� ������O�f�E ,�LF,oJE��5��d�H�r���/��b~�&[��A�[69sޭ�{u����\ ��k\lR�?����V2�߮g�YI{ͽ<fn�T:�������@N�ɤhy�����ɖ1���Ťd�H�I2�]�+��r�-������M�'��g@���R�s��=g�)*���R2���ƥ�tW��ïx˦	�o���@ʫ��n� x��k ��rq_�Ʀ�5�"�z�I��0�I��X?�0��-I4���@���Y�;N �����������d��_`g"? ~��\=�����M��3��P��X�����z.D��8����@0��L�cll]�����gJ޸���w��6�����vR�!���y����X/��K�a��A���G[V�)�Kr����P�T<�{oU���?K^�s�FWivP	:�yK��i<��M�G.�AC��  �Ð���Yo4q �H���[����E�jɁ�F��|W��;"��*/8P�|�ԋ���灴ֲ�/��o<Ʀjܝ�¨N�k��C�~j	LBRm�����1N�ԣ���	4g9]Z�������4����3R���<V���%t5���ë[�������D0n�ɿ�p}�4�)i����/˟�5���V��7%��m�dS3][��osX�*{�PJs`[3��{$쐽�粰q����x�?F��w�`�{�O�<���9V�w�ն�~�@��n��{qk�LQH5���<k���,�c׾�,��� ��|�g��]+c���44�*��{%-�\���	���k�Tn��#����M��TB$ W����rc�EEљgA��r�JAP*�n��5g�3����s[�	�!�������0�����
�?��
�U�]�b�DTlo������TFh�0�AC����00���E0�5�`��;]5�&Z����P(0/ w��\I��k�,�������ߓN�����8	�76�@�QXC<�o����:.�b��pM.�{쏩ۇI}�<c�JX�;k�����!ď�=s1���������#�b�CH�W5c�����#��w񝯜�H"(L=+"ea<
�c���\��;� N��hE�!��1�����S�ߗ~�<�����ZP�h�ق4���a~�E��+BE'��^�B�^�ÌeP��z��U@�R[��_ݚ���9n.�YEj]��BY�N-�L���t�t�j^�2�W���daec���z\�uzO��1x���k���>��w��&o���^c���L�/>�O� �hv�����f��oX�H�Q�	\��(�|I]�I��npmEh�C�{�_ֵh���Xl���őר�xq/���)���Ñ�}e*�f���]��m����59��	���M�t�@���%��2X����p@�K���}�\�����24�ߓ}��t�톕�������G�Ý��E�����p'&��}�C[����Tj���gm
��U㱣�RQ�}2Qk��1\C��N"�*Ǘ��Q����������4�6��%�zy��RV���U�Q;?$�*�Vʤ��e��0]�m[�hv)BY��s�zxb����%�\��(R�y�3��������]U�枻�a���R�\*k��"�U6��7a��s��&�>�9w�Ab�<�v��ƀ�����d�m	�>�n0�Ȩ�X�~�D�h� ��6Y���>���|�~�ѓ*g8!v�$_�J��+%L#��vC-�y5���r	P�rC>>��7�w#�P[��:�=(�Q�=��i��&f�??"�Ѽɖ�6ջ+����ӧ ��-��T��US�~:��o����
�� �g]�d�SL�7��o��ߝ�BXmϯ�}��9o3�<�[V�+\JM���Nj�.��|��d�/������ �俛�e`�)2�� p[T�-k����ި�_U�2�~X��+�*��,q�a�����wa}��Ć�u\���e�W���&X������aA��>fH �E��6%�9��.2�u��a�g=�"�p(:慳�k��Јʏ�ι�4�~B��٢�+�������Uy5y ����PQZ�(R.E��n���Ҩd�mQ2�lܰ��u�!mJ��7�fk���	�����Ps�P��ɂ�|�&�%�Ƌ݆�K:��ШpF}s�"뗂�q}��wlؔ@�����8n;�ʬ�O����x$Q*�=ҕ-�� wcj"��R#~�$����YY|g7�?�=�����bφ'ȩ����4�T�mS��w�P���3n]
�3�����/����fZ��egnUUVa/%Yn�Y�m,-g0⸗����y�Ё+����ѣ��>�� G��o����������ᙠ����3���{���B%�)[#��\i��M;�JQ�AӍ!(K���vt��X$�׃�-5hu��uк��h���o�`BPL��/���[���V�ͩ�/,D�1B��L"4=��տ���S,�
����N0����*e��{��g�sK�H��L::���k��(P�-�B�4W1�6��e��M�>W�z�=���w �^ϡηkF��x�B^*�}���.�p�8d�W��;��2;���-f�ZB��q���ݘ��u�z-\v�]�=�Ya�4e�M2�*��D�l�X�Khڵksm[2����v�ݦCxHCzt�� ��
b(�`�%ρ�F'8��Tg�]��H��~D��R����9̓���%��=ť�=&���.��[��OM����7�X�,��R�C��x�����zp�����/Eˢ�/�����3VGSj�,`-���|N�:&�Y�_cN�� '��^;���Y`a=b� 6�>��"`߯�Öq�5��	Y1�ZuD�5���|�� ��:{���v҂Vf���r��h�yh
(�l�~����	��c�����-V/$k�C��F*��u���E�^�YD����M/o��\`:����.�.����)�j�.��j�kC��+���G�_Y�.'��h~`���c*������Ъ�Z/H%  �ҮI��퓚����������WO����Fv5/9�����{�>ZXj�����od�����k>@�M�KA#�ѡB�Հo�+����ƕ�>���8� ����S�	 ���4$y���ci��]����W4-��H����5_>}Գ��Q����d�,l-��j���������l�ݜ+M�Ҿ�ms����qBM��y����>���y��\8�V�<<�~Ns؊��1̗meE���w��f͗�B�ċ��.,�O��헙�w��`��v�zEN6H����*�#���k�ߛ��/=�&ؓa�x���2b{��I�P���{颱��fC\���HH4m���C��L�w��k���ߕ�y�������c�YdMϞ���j����l�6��ݑ�κ^M��6�Ǫ�~����!Y�+�-C���e �dn��l�@��٩�p�6������WJw�j�.� ꮁ�c��X /M�x������-1���4�Ҵ�H���_�@�H��a�Jse�׫&{�4�2��"+�~�۷S���hpdP���j��u�H`[\5�Κ��k"Z����$�����/e�yV`�Ŗ�H)���J&�ն����HO��1Yq�K� �l�'��up�q`'?��`MpG���C������u@6 �<�M��o�i�M���;���S����P�����v�Q�5�ˮ0�Y:M���u!C�����E �+sy7h)ȃ�/ 2HR&S����F���rbڪ���:i�d�������W>0�����;��X�{)���A�:��d�Z��`V䚐�Ο�B��؞�x�,����K珽�� ����v�>a�摯j;�d�rZU-}�uӜY���[Ysqۉ��=-�ݴ��d.���
r���!�pi	Dz�8�	�眓�ٳ�Z�{�eBy���O5D��.�!c�����8��o�H��sW�C��x��Yyny ,!<YZ�8��Ł+!-譾��U�$�Y.���a�}�L�*�'YW����kg<�56aV�ǿPlװV8�s��*��="���?�=-B9�-�nx� �(ۛ5\��w-��2T�?� �Z���fj��
m�Y���A��X+�;GO�%7q�[�SO[�vXe3ׂ0I�5�}Zt$�1]�G��
 5��,���t`�����Ν^�Kg���. >0��]f�^r�*�Sj��<�+w������+�E�ӷ��}���~p'�s�,�J����)�|�{O��U���ߥ�G����:F�5��ɛ6�҅���p`٤/��řk9q�e�8�L#��A�3�g�H�Hyy��b�ǯ�<C͓ �dw�!�b���z��� )�nXb��%���%Cb؁ñ�����!L�p�S7Y�;S����n�6�+k��?�``Z���vx�X���W1eҨ��T���SP���;�S��#l�h����}Mk�@a�F��Ol?HE�6n��-���8�Ɣ� +Z����VƩ�
ӜVw��>�q�k�N���H%���U�{�J�i}6Cb�8c�����!����j]����@I�~�D8׷}�ǽ���*���l>�"����R������U\l�D�Ȗ����o����)�p�\��顓�㕕��(5�u��aiᵾ�2��(��P�E�&��.\��3����?4�+�W"<�5��'!�?�(�e}���f�.�e�����_6��b�݋�>�efڂ�T�Fu-Q�A5i�{��A6������׭���Vtǆ_������n,~��P:�wY�����]������x5\�k���C�:nVf>&��QVQ�o�{[�� ��9���Ծ�8eI i�n]`%��A�/��Hڱ^�,��g0eWr��O�w��^SlJ_S�����Π����2���63�=WU��p��N��>[Ɯm�ƭ�fn?�օ��^E܎g�m���WGr6SB���Z�/՘q�6SX�[�ɀE�vh�����P �{x��_n�s���
U0�z�I�ø�8��B5��B�dE����5�ú]ڇ�w�������^m||5+�{,{3�v����v�F	y��~��Lȋ�A˘�z
+5I�! �kI�絾�%���r�����}��o�3/c璁�
b���M&���k9{��gV��\57:Ɣpz"�Q#51N���K$�,��{9W��rLܴ����^a{�P68��&��Z�m�>︋�[K 6��̛���h�"�-2��n������`�EX�Aׇq]�	b�ݰ���y/��.@TZ[o��.J�f`?���yLćo��L}�6i�����o�νSс���!nT�QYٲ}� ��Rs4q�b����ʫ��7�=�����S���J���wi�),޳�����>y{���ꔨ�a�S`߳���?P6=��㯊����T4`3�t;���A�fC�*O�d�����+�S�1��I�(w�璧JQ"?64c�<��񑵆P׍�V�����	,/�3�C�7����	2\� ��p�����e�-�'����5¢Na��<�.$s��6-X����r�V�,�.`����e�T��TM�C���vx"���=#�3>Jf�;,���QH�����;���Ŕ��n.-՝��b�H���-��	۾�[%�����Pw�l	��5_�!\-N���� z���������4�%_+�iH�B�X�E�BcV�����@�ӏ���\^?ߕ5_l!�9��
�U.��6�J 8�N&,�7
��KU���};�jLYg���
��bPmփ�����J}�)92�O�-t���-���Z?������h3r�խ�Cj�ȉ1�g<4�%�*_%LVm��t�I�d�U{wq���G[-N�(�6١5p�P��Z�GB�N��D�1Yh�Q���Sg:�}	߶��Sz/�ҥ��{�5zU�-�^ߞ�XO�bp;���������)i����=��'�͊|��2#��ֳֹx �����Q��Y�u��`��[5�G]B���"��:FU�nb�أ���ű6��~��:51e/J(�$��2/݆'g>?H�M��u=���$J�ǜ�@Z���:[�$�f�42�{=0�	q���p�{��s/�Uu��G��K)7'K5$�}椩V?������h�.
�X�aA���R\ը�/H^� Hq�th�@o��IN��t=��G#6w���}���YZ �z�,��?��X�%+�Qd�f^BsVL3B+����,�jF�)c/�t�ͼo��7�z�ǋ\T5��^��m�(�#��"��8,��೑=y�}��H�#+�*Bp��m�L�5pR	r���D�Tj��1��		QO�&�?%3����wB�7S�RK(��g�t�y7�d�d��E���P (��-���5���~���Ĩ�(��c�MM���t�3��""��0lrּ�ր��2��힀�O~,]�L=LN��c��H��I�z��i��r�0I@��C���mi�M�I�<!��	&��k�z7.�2��#Vw���ۮƊ�"�6A#������z�U���o�Ƭ�:J�C�M��0ͨ�{����;9J=[Fp�V�R},=hg��0�� $�:�FWgYx}Ŷ�W�';���R�����{��۝��w��Av#)l-�|����]�C�jM$������#h�x�胤���ELtl�}?+��劐�>a79�,@hIG�)Fk�:�nX�\4m_��l�~������~{�	��F'?Ś�/�9\�)k�֒7G�!zӍ*Ui����6,�DA�\A�Pz�k-�/���������9[��]>��Ǒsk����wo:��Ê��ّ2��Ⱦ&0H�����ũ����2�0��0v��3�B'X'�=
Y��	�o����2�/����˯Upu�n��7�̤%�yP���N$��  �^�bc�� ]���9zH�c w]M5Ti��G�!�+�*��Kg�D�(��+���F�x�+&�����3+'v}�ifl�����Am�Nf]!+"�湄�&�-��P*�1��q��`s�餱W��6�p�0�V�M)ĳN��:^�^�[�\���7<F2 ��3���!hQz�b��M �>+Ɗ��Y�_�ǳF��"��EL�������c����T�H�m�<�'������JLR���>WMq;��$%�D��$��C�z�s[������,f!���M(BF;p>E��m�w;�j���wfW�^Z}���Cx�&o#	A� �1�m��o��~�f��_��4���
a�P{f�vKk7K2\�l����@�:[�S�E�dm`�+nY#+��-I��%�t�S�C������w\5d�]���c%��d��4����j�C�S
{X��4�x�,��}�d��{3���=����������L
}�E�+�e�Q(�F�30\5��N�r۰��V�O�x�ȼDG��!�q^$>� ��V���#�Iz)��tQ��BtI���aӽ!�P�������2��K��?��C����oX;>oN�Uٸ�~ �)9p/wL��	�iA���6v�lW�N/�d�R0��*��!]�^1�>ٖ?Z��7�U�)�s��F�%��x&���D��<���^7_����G� S������[��#P[6�<�[����2K`8��D�jSHZ�3Q��RV��� �}����ar�}�-�z�t-�/=7(�������E�w_Z(�Y����l��5뒆Y�S"��C�]V��F`ď�5���@�O*���m��s�;���Ĵ��	�����(8Y'����>����%Ӓ��t+"b��n<��A>o0b��c���?>t������y�fף��Oi�޼�%�Z�nC�߃}�R�`}�|7���#8��ׄ�Y��;7�V*�XWa7K����LhJ�C�G���2�UT��_g�G�n�5��$|!�GaW��Tə����l�#���=hQ�V�~�<"�~+ݵ:���w14��G�%�l�0�I˜c�Z=�D�As%b�x�q�ݘN�����=�d�ԙ`��Y�q�[5p��ÿ�P�e.�����j/.��#�C��z:��/7/#�G�����ͭ�Dᠱ\�M��ytDK����9�)� ����@e�������4���K�=��s�:[5�zQ#5��ּ� 3���C�Zul�ElR[��l,N+��U>����c��V>$��9@�1�U\��F���Ϸ��4�N���-'A��&����J*+xM�_X �ϡZ	��{��9��yJ��Y:�҃�v߇B2^]�nH��i4���ߩI����_
�@��k2����A.H��ْ����J:��X��ٝu��4*��`˂NQ��lc�Fn�5E3&`r���7``8N;�g�����p�uh�g�z�g.s֮Y*+)�O�#�<�G�%.Z���|2��nbF�ݻG̲'��%R	>�����2��+�3*˼5zw%�y��B��y�$�����U��y�q��m>&�5Sh��q�.��l�z��O�!�!�=)����D;���A�C�5�ub���u>"���v�`s�����G��Xwf��/ĵۋ�0p��0d�qD��N�d�� <�ni��6����W����^�����
;wC��_#�!��@ ��=7��F���c��g���y�`���c�!��P/�o�F
!�"ʡ�٣�̸�u�G�d�U���T��}G��E�,ď�qZIX�+�H�C��7aVq3b�q?�Hg%����VM@&f���5�XM��ws���SJ�t76G�����c� ��]xPpH�i4��qR�R`+�!��@�(*�3>Y�ZL�~t�������lC��r�Jv��A����Ԥw�M���iKl-uz��[��@L���!��Dg�a-�Z")6�����;诺g��N� _D ME�<ۅ�,^_�nV$��7-c���s�-�E ��i�\xM��]e}�-�#�<��E\�m�����J�6; *W�a��6]�����	}|���seE��U�+V�F��:A�|�_ҿ�� �����^��E���28
�[���[�E:4̡�Y�'��Y�R��1L�>î� !��'y8�e6(�h��K�xG��4Z��̽a��H5vPr�0)D�Va�5>���bJ�VyKݬ��A]��C����ǣ48�z�Q����QnP
����YăG�-�ELɁ���2a�v�������8V`P��f���Ѣiz�����f���hR혰���������7�X���x�Ҥq] i�i��)3q�v%�6ȊĸUvYt;g0M�}=���?r�" �:�zg� }'?W^q.�e;1�����:U��J��*,��i����N��,���<�xB#q�[�����1@ȑ�I�?���*F�ڝ9��A9�jpn.i}f1aYY�=� �׌�wO�<%��m��9{���'j��L�`�R[�����3��0�����R����/��_�w�m�}Ɨ�T�4I��0"�
�.��&���'�f.I��Zw����(.����q{�/1aMk������.{��H�����s�ml��[�8��cYŐ�N�!8��tե��;Ȃ6EJ��mt��mW�dER�zG�A(����mL�u�+'�r�A�W/u�B�����6e��묶�r��eBj���4.���ø�In�ֶ�Y�,>*UJp��ȍ���Ip�+
��������.oFZ��� ��W���Fh��(-ӟ��O�Z�(���6-�ɴ2��1�
52�~ز��Do�T&�a�0��D[�k�=ʣ�����B�`A�����ɌyN�S���þ�T�Uҹ2X�ה���e���/��.�v�jm��tٴb�h���٥G��!j�R5�}��pQ��]1UM�&��%5���K5hg��f�#�]k������-���T�ax5�dB��o���?!� \-}����x��H�%����{�S��h(L����J���<ɣ>��Dzp
� Ds׻�%�ˈm�q�"E�0��b�1Z�q�G�e�7I��:�`�
5��`�ߞdkҳ|&�r|����>pL�+g�/����^�R�҂�1�̧r�(�Cn$oN�0���<�F����I����zF[��K���}q���t�����#���*I�B�!�<����f[�2��d���/<B%J�l�A�n��a�v�q.:[��O�k*X�N�u�h1[B��2��N�N���g�u�M�A%6%�8y��a�1w����I2����!��Q �Gv����fd+M�1Q��:DPвLnY�@��ǲkk*Yy�mƉP�	2t9��(PA&�{(�׼�;��!ɨ-5\�)�%�O�x�%�AL���mm�F���'���+e�&굶GFFB�{uO����Qc�)t�5!|?�U��� �a��9� ����vJՉ�7;[R�A�E�T�CE�N|ӊ�����l����nŋxTT��z �;<�5��hn���t���� =dr�-_�zHS���0 �*�Th]��t�c�DnnRq5���ٲ@�����Y����ǃ�������#±ZQ�n�O�/4���������
��5H��e.�p��h�C���<���T��R��M�P�@�sAv}���ڲ 2E�d�c����V��4)�1�a&@�m�qT�[o��JH4���� �i?&��],�J�:H�����#_	w<3~N˛9h7x4}�:�/L�O&�=KLy�s�T ���\�N���N坳�Ը��#����`�}�g���9�s�5eT�3ﴈ�����X��t���'����Zx��G�}OU]�x��d���2��"�|ء �x ��pv��w�Z%!f����D��e�+�E�Jcr������^k.%$��t@Jv���l ��,j׆(����cW�As{����o��V�E�h=��N�n�d��DC=BS'���
j&'��[09j�����T�����G��W�1�j�����Zf_5|{޶=E2IX��xQ��A�8"7DHW��s,Lqݿ�!� �`�Ok�r-���d�7Y��	�)��uk�P ��(;yZ�+k�i`�������/#g�p}������}��P���*p��N���±IF�h~P�Q*ǧ�	`pJ\/
��F������:�=#F���5��=[�\x^��\_�_�ٞwQPy���Y{j�H�:Kݷ⇉�$a�/I�q�x&���z4�( �-9�ee|��ت,��k43Ѥ��DJ��D�]���-�@�+�Ñ�ZM���I lԨ����
� !��Z�?7|�/X?�8����B�YA=�5�3��lK_��k&%{�M��SS-ֺ���X�UQ��B�j��	B�I�#��m\���+E�����=J]��-yB��J���6�|xm�`��)�����K"�4f-m�|'��s���c�p�+mAۻ��ݍ���b�4h��V��.P'��'������ǭ��]�.�P��
r˿����x�F����V������d��ڏT%�����)L���56*��a&nQ�x~�(�^�6a���yL�Kz�d��㢯�
Rt��������Ks�����I��b�{I��ﹺЁ��{g�4��İas�p��g'zb�Von-.���9j�
5��+8�O���NС�P	��}]�Wt�UHɲ�3W�=0���ި|��G{���an9�g���%SlM�G;mS4q���y�N���oӭ�@�6ݐ�Q̕V�_V��xx3�l��<R�.��.��9�茖Z�b��c�>s�i�[˙�t��#� �>N��!h�#�|����d�=�vmp��~��v��Qo+���`���v��*C�)S�i�����?,g����7�Ȑቿ��L�A�N�ݷs�2��N��
��j���SQ��N���4�=�(���w#e��&��O�� ��YT"_!ޡ�*�)4[�w�8�\W������*��� K�9���#�?�Z��ah�q~��ީ�	8}�Gj� dՊ�z7U�8��"�i1�(΢l�L�Z�/ȭcRu�h=�����5]��l���\M\�������6�D��9��`��G��D$�U�2�(`lz�I𚞃%�%�h+Λ�3N
C�N�Υ��
�3�����|�Bx��s0�rGO�zlT���Y9eK�A5�iY��F���y:���A��N|D 3k~�R��L���΄�WǵfҦp���ȿ���"�@�E�޴�O3pL���i����5�Wb�_Y��ޏl��N9:p�I����$s��4��58o�G���O}�����2��[9����I,���mp����k�e������;U�^���%&�+E���y�g��d�)�1�ܕ��[ ���	��L.�=2����Pkΰ�avuv�<^�rZ�\�02:v�s�,)H0���~�V^`c��u��ժ�̙�IսQ3�Z��XV�b�c�'�VT*D�w.5�5n����g%�˓���:/��A���}�P�Z?�y����Ѩf���U�� sͮ����ymB�HuxT��8nL���:��?� M�$�ÅJEd���>a{�����!�x�ߦ?�D��V0c�[Z��i;1yG(�7�H�|m�"}���}��fC*>��>�ҥY������$	{����-+�" �,�I}�ua���$gf���	'VG����-���0�G��2<%��.�0� m��!��J�E�~��L'�Ï��S�gс��'�g���M5��vH9��mG���4j�E^ΠF���-�VΚ�K�ɞV=�,3!��W#�5a�׋xLtzN��R��G��P��(���P��X����(�c+���he�,n�[��:�@� ����2GK�^��z��a����`BV.Oh� J����J����2�ђ��;�$���u0�L\5�W�$�/���@�`?�Ļ�oXq)���8^�ff��<��}A��}��b�|~�5p�V�3� ��C-E0�o
l75XN��TD2�)�zOu��5���K�ǆ.Kz�Zes(�L����-��"F��=S_wGk7�f�6�e�Rt	�w��h���8�$|؋H��/��)9N� %+�6$t/��.�D&L|����Z%9���(�ԲxV�bɫ��l@�$5F-�[��V������3����{�y���0�h֒M������ֵ�2���*mX��<�o�7szq�~tG�w�B�X��?����� ���C���L��6X�r�|�O��vo�C4
Y�3p}.��3.��EB:2���Sd���Xkmpڬ���+����y�'R�d稽�P#�IƐX�b����[1�UuLH�tIۜH�`��C/w:�1��<w��v�]�������08@	���Bz<G� �[������y�K�	)�����nZ(�K��48��'��26��	{7TP|�ͫ�27A��D3��mÙ�Y���M6�ڪ9�J������H�*��{�tf��CB�9���t�=^�HAG��]P?F0�c�A0<��^"�|Y�y7���]����:�.o�0���9�U�ڷ�d0#9�A�d�_@U���� ���	���߲�b�ߎ�4�D��;Fe��c� #|���j�GP����l�Ԕ�3l����:�k����B)��%���̷�o$�mDk�׍',��v�	����/T�dLxn�m%�C��a{���U/`�����=��x<��:���ݴ��W����ya�uS�*p��V�������*���Q��:9Ӂ;5|<��P��D�s�'�#y�A��S&N�@1��2@
��q:��zS�@"C�1�����c�u�����̱�4k��o�^K�#��Kxp۱kZ�_N��ѡg�]�"-D��It+o��8X�-��Y�lW��(D1�M�v ��R��$qK�<UP���Vy��;�n��@�V|� e��:�z(�xP�͠�;~.�ت殬m�d��gg`�*�`X�_��7�B3�i�k��K��]'d�?��'_+R�p������:����-#X��E��
�FY� ;��ɕ��H�a)"��-�%�0���Q�Z۶u[ߟ]��rQ �*_D�����>�S��]�A)������<��'�<GI��4���{ ZBv���<�����/Y�]L�	NM��}{�ūkׂjF���z.~��\������puo�ᯚ�T �/1ea��1�,*Ɲ��K�Ok���g�=h �'�J�!�=Oy{�u���&bf ���L�����N���,Y����k}4͋����x<��J_�$`�y�m
��}���⫥�{��Nh�7�~`��V��z�L?A�4b�4M(ȚV��59T����؄6�f��φY��W`���1��q���TD?���r�n����Ȃ��ܹ㳭9��@Y�9�*�f9o~�����ٷ\K�H�H(A� *�6����w����*©���Rv�;�9|w�{�W8{S��������䊪B3t��NOTq��@���ҽ'�D詠��|t:ȧ�c�-�id8��t��d�ώ6�T3\e��k�cMT�΍e��'ۭ��X{�����r +�i紦�!���f�/<��9��uo#KӪ�Nj�u䷐G�Q!j)@bu��*���Ry��yG���H�F<�ꏴ�;��b2�(�{�Re�5����)� @py���2��hȇ1��5@j�ٯw�u^�b!�ܭ���E�+@Rk���x�n�؝|�{��-9�H՚�B���$��w0\gB9��!7	�nޅj��$�#����^�!P�<n{|[c�3|��G&����`9t�6<%e�+�h��E��[!5`=�e�0�����03��q��O�%GP(|z��l�MX߭��Ck�v՗�� s��ʬ�.�a�E��l�prG�#�w<�I�'Q���T�e��Ͱ�sl�M��t?�.4��,��1f�
�`�ܸ�-�S�=�n:�~Nq��{��M6s4軝��e��cf� YV�Mp�ϯ��� ��C�����!s��/�	�͈��>��_l؀��3��#P8�e5m:r�\������9��m���]��I�D��=c�bI6u.�Qjɨ��nݜ�U�E��D�j�m�RlD�mc?|F��O�Mpo��S�/����ZZ�&����q:�c[�@M}cw�����$jJ\�~b�`��͵�⾆�;G]���(��:��>f�����eSa-�Kk�Nk_p[˒n�����IE�5���,�hL7zZ`GU�ޭ�l>����w�)�p}�(��)���BD��x���g� A��
33��U=�@�R�#0��W�����N�j���	<}U`l����w]��)�F�
��/� ���WG.��޻4U	ڷh���r����{��<.j��w�ʜ�Q"��p��$����@L8DҨ���ᛌ�e���kc�{��|*u
��Tj�V_@�l��o?ǕF���0;8 T�Y��c��9~Lj�o�,����A�c,�3���!�mCD<�#�ˣ�Zɪ�f�S�f\��B�V,3���x#����4��>����S��2h����R��#��Є�<;�\�L��δ�y^wx� `�����L�g�v����.._YW����`���	$�d�*�o&��?���0�����h�i�v׏9]D�����F���O�c��?q��s~��W�ƚtMdK3$����Q���8�"b���Z����j�L4��;G�-X��AK���l�(pnA^���]�P�+����G��u]�X�)���
�e����'л����N�����Ϝ0>�B�<��ձ�U��n>�ljB��P�<�N�l&A��D��Ԣՙ��G=v��hc�{b��\/���etǴ��-s��.��A�7Ŕ΋�a2�#�7�g�K��u{�"a���'Y�מ��Myr���-�?�4M���@�RA���/��եF�3�gj�r�u�k������t��/�����<�C^��a7�U|>Jm�$@���n-,�ד�u���J�,gMnR�:������,���ٹq����-3>r.ӵ\�p^�B�M������*)�Cv-gj����0f�X���i��Y��>B�X��D�ۿ�l'6�h�Pt�Ea��\&��0S���3(����D��~��^� Y,ѓKV���{��$�R�& ǚ&�gܹ�ˏ�)X�ըK{�J��?�l2K�d&������B��)z�>��ng�H�5�9���&;F�t�� �-���`$����2 <[�1J���4���e�:���9���h2����(�vY=�:N���tE*����G@OE7��p0�E؊��x�y)�Fe����{�~����U�@��Q�6�1Oo��;|���G�(���(D-�Nb����m��ϹNi�yb���~~���\j|kJ��!o��[�IM�;H�E�U���u���H'�BF�L<��O��,��=^�ъSH�_U�B�e��5��b�ILU���&.W��e%�p���(�ؙ��L�;ܷr�$l���{�i��v�2A��2��Z�O%�����9��\=/i�f��翊54|\�ss����d�6+1�0�e8�|�j�,�G��b�W|3�mZ%c�g��J��"���H\�m
���0
�00�+%�HL�r��}����w��񝀼�%@���ܷk�����9U���(�HOd��~�7O�89ټF�$��H��`?ǘ5�kz��1ם�� h�;\�Է�M[��	b3����*�ˆ�\�	�<c&�!��U�S��a�.�rJ��j-�t/������Pt7=1������{K�x&�={jd E��[EЯF'�0l6C��N��n%�#��5RrZ��+�Ӓ2�(�֘��W���Dm���
�]�������l��:L:#0ꁡ���3�W�^pDA��e���롇Z�r54b� گm2 Q�����ԍ���jAJ3��l��O�7[�z�C#����<�,9
����'��A�����_�EBr�i��b�L,��PB {�]���n�{�2ty�� W�Z���S��p���q{XW1?u�I�3�h��	���`�Մ%Ɣ4G�S��⁄p7��?_zb(�� =8G��3�	3��a[���4�,L76&SS+�ݢ�ۘ�i,ҏ+����j�M��@�s�ܰ�)&)���h:�+���/+����N�Q��7��hb�4�jy�ҤC'���SW�U>iR�D7H3�t���2�O:�ZD��}!+2�_��4���S_c#>ek�c}ܓ������^Si� 1	�p���0	'S
��}��脧(J�G$�I��$��[�ٹ���⒝�<ݘԼ����#��?��:�T�m�j�p��W����Õ�lxIΖ��~*�>�O����=B�MT�X]���n�ߙ�;��й�Z-��M>�s�Si�{��7e�����{�(��#7i�Ĺ<�5|M����֧�^����1Y	8�C��vx/tĘU�?L=�,�BB��;�Ěo�	nf�#/�M�r�u�ǰP�V�8�]���*�֦���/�����f��q�A�P�Ҿ������I5Xq��.��6�HfNY��
�G�Ⱥ-�E�������eV�R�N��c��2>cв^�����$�G�|�u��4A.�3�:R3@�fW�6$�G�gu4dr����_��a�K�|�S�Z��sYk�}Im~;��O��B+2�#0,�0 ��'/�Qؗ�������U��r�K�q�:?^O�XZp���ƪ�6��z�$��� ׶��TAY��@��^*zN��03s����JBbی���F�z�-ux?�"�+~�$3�2�����y|��%7֧�>��a�8p��h�#��c�=����ô�G4+4֠�J6�kgL6
Ni:1�I���N���0~�8�?L>�($��Ѝ�X���u���s>�q������, _v��2��}��s���M6��z��@ �V�+�*�}�Z48~�0x���;��BѲ�5H��r~֓ V��m���?��BT1�Bw��Y.�D�Wh ���N �a�/�6�p�0�!~ѵ��@�.��S��nf&��gG;�0�,)"N�t�U�/4X$F�if�#���ސN�I���q�ڔb��e���I���l�ep�*����Ct�@�z��b�%��T��'v~���c^�r�7Ry�k��B�<�tF
;��#���`�>W��F`��@dA���2��XB�~s؀&�Q�v��9�0jQ'�M�7�h %��k}��E,Y����@�����4n���VL�b
#+]��	qL��j�7��F� �)�"�i�k͒S��i"�9�;��K0S����+L�l�uE�%�-�R��k���{�c��# N�4V���z��R	"��4b�|-UTM�L �v�� �;Y�-@��?�I�+��r��ܩ�B���������0�6��9 b�ɮ�z���c=a�d�T��jz�������Os8��;�<��x�>��O�ͬղp��T�O�!f�������IS�V�Q�)h�_����P�U�~���,����S�{Qw�5���[G��1����z�.@}���ٲ���{"���\�MNCD��o��ԇ�W�T�.Xj#�mbǍ��T�A����Y���|9�q��$�������	���[L�R���EC�eE��|E����o2$�����F�E�޺,�тy\��ɞ�`Ezr��>�}���P����1v���L��0Z~`�v���|��N&�������a9��9UU�F�i:0��Ƚ�V@�7�W!����B�ꦓ`�A��.Ŵ��rZ<h[bǳ�c>]νG6S7P��bC�������Ip��nJ�l�!h��NP�-^�x��{~Pm�B�TS�W ��P��+>�FѶ���+)�¶���+e��o�e�"%��ִ�/�m��̯Y�G܍�t������Yd�X�'��HE��ڨ�c�؋b���a�$���`�^E���{�F��%�[�_JJHesTPlwl;w=��8�O�2θ�3��N��]��}��+,v[�X����'K�.���R�0'
I�n�B6��i��~�*.���2�oE?*k���J���_�<�ǭl��Oi�/rţ#5�G��W��IA v��[�ߔ�!�.�^e�%7�[�4�Ie�!���&љ� @���a��^"o�;�k6����eL��=�	�{��eE�uкΉ�u�T�3!I�C�7�r_�K;Ǥ��663藞��_��;e�W��bMX�dYg_����
=��)���
����Q𸡷�Bl�~Iuk���XH똂^A؇B�"����C�r2I�zj
E(�����V,h� T9��1����`JX�hG�hM��R
's��Źg���~s(I��N�Yv���!w�q[k�
�'<�;ѷt��K�I�..Q"��=�6�=v1���l'x��D�%��)�|�%6:�%��|����`��ǹT�,RV��I�EY�*p>���M0�Tܸ�wm�Qg�p����[��p�%�#�o#X�������q�0�
 8�8���-K*y�PΒ^�=bkg��7�a�
���7����
He���E6��o�TrL�˲ ��L�-�����f֊>Rmi�g���*�A�>�`�8����Z�Yk`��༱�r�il�;�K�h��yG偸�A�w���Ѓ�(�'�h���u�Y�kſ0��t'�1%�S*\�n�5��oq��y&I�>���8������.6h^�v�j[D@�4�ѐ=H�o&2Q�!յ�"]�;"*�aG��n�P�tu<��i>��=�b_�� h�|�)��[
�
��D��>�ee����ʹ���:�ԔR�m>�:�hM����;X�gt�"���-��12/��H����ΩF ���J]s�&]A~־��cZB����MT��3�-K4 �6�SS��[�����}	�Dg�pO�}�� oL���[��(�0��.�����G#�E8��L��R���mr>��1� !�t�/g����x����f��CL��?T����Or�!�a댶�JLC���nn[����KCm�_/��"�W���`fأ3ݥ"�3"��_��*�|�k�4VNb�D'H��#܀1�d��^�� v�@�,\�F�2��邔��3"��نGo҆������Ӕ�/�0���v�_��؏v!�5�,ƝF���fVp�ʚ�Ό��\3(S~��vX2ϞT��j<�ύ����r���e\���"�M�:�4cV*}�rb��aY2�cq�C�c�B\���W��`��Ă̘���UZ���VȆ(�������l�d��I����;&XW��)O/B'�:�����e�pF�u�D�M9��P�s�!�<$��w��j��8�aL|�;�Ĕ��`�CI�j͓�FR}�jEA�0x��(J�!g�<�B�(�u4mI�c��Q�8�J����g��O
�9�0x s���<2ը�+�"��G��m �f����p�p�{�_u�,��s���W���$𘳪K�l�eg��bҦ��k�m��`p!g�D �[
nf��ͳc�������ّ}ψ s���@ŦM��>f�}Y;p*[t�/Ċo�l�/fڵ�6tX�e��/�b)�4��Usϩw�!�Z���繳���,�5K1M**���g� ��]�:h�'�ӝ�&Ab�DW����"�O�� �W�0�7�v��u6x�H� s��E�h�'���wlǟ�l5y����E��>S����O��eG����ʚ�"�t��Q�LZ=`��RƘ�M@�z&�X��'���r #����_o2��Kd�˝�}\5�������͗Ռ�I�W���|"w����@�7�>*1(�*�'�����cq)lv)���M� O���B���pOHY��b�b��@F� p���i$����W����?{�3--�m���7��wA��&Vq��7`԰��r�*&��씢�q/�B��O)J���UI�Ձ씆�uG-$���Y�nE'���BC��[֣�{%�l٘��\��4~�[Њٲ_T ���{�;���b�Z�����h��<ccqqƜ�1<� �~�l��5vo>i�lR�xś	�\����kN[eլ�S����ujq	�T[�3Ӹ#��Z{��Z8��UT�J�Tܪ}ȣcOd���Nկ#�F��s=��}�&ll�T�ȉ�����8�\�ޥ��ܟ�9qm�Gi�2�N�)KMNl2}���r�Ah���5�Ȳ�Xe%w.:
4�$���|��Q�f3Ս��Ѡ[�` ��iԻ�#D����A��'A�]�?�����<-���e]68g.�u.
$�a�/f��-A���a��BK����V��!C�.q=;���u25Z�HElX탔\Ԃ���j��+`>�0q��b������r6�>���tW����+�`h�v��9��"5���DEk)���Q����*M]�Åd����S�c�f�N��4���
�'�o\�P�GB�hCm����ޣ���K�4`{�H6���D�#v��y��}��<�5%��Oklx��kQBdf�]�B�����K�)��Z�p�J����j$�!�ƥ�Uu��O?F��V��t�+��w�ɶ�k��#@k)��3��A+)~��s���	�M�v�����-af��mΗ8���3ǟ�C�e��.�or�2dնm�0w�O��P ]�:�_���QdM�Cp���	���o���G�A�h�Q��v�]�S��z���/�m�R	�_�x��{m�;�+ꔙ3�1��j�������0����9oR����aW��!��ٜO��g�.�H�������e�&���D>�JD3�9��З��u���Щ�Qح�v|�� _!����V#s�ܔa�\A�������^�wl�}Duu}�в�L����k̥�Zhȑ��l�N|���gA��x����k@�m��G��p����.��7�?�u�m��/��Ιݮ&��_hQ#��:d͈d�B�	����-]�.��3a30��$YiEE����͒�4�ɫ� �+� )]`fw���VW�ڐ���k6]�e0� ,�^��>"�%�7*_���T+)�ٍ������u����ǩ���R���i3a��t�L�)'�;>yd4�e�B&��aC�1��ʮeu����w�1����}=Z�	�_hW���EM�pU�	=����U���D��c���<f�'Qh�cƶ�6řjD&l(��1��kꗺ.��RA�fĶ=���؊V,��� %�3�=��x���0I�'C[��Xk��Q9�i��"|��_�G�-BF8J��e��J��bo+��~��ٓb�t6�����.����b k浶���ޝ��,Abl�h)xܸ�eel*����3�o�qAU�3�5�>0ќ��+~B����,���ǌ�Tu3t��e��><�k\PKUV}B_u�kKI�I�H��SL�X�x�.�\O#97�gb�:��]���
��� vC�%2����%�h�'d�׶CD�$���HUՙݗ��J���l�]�{�8M(��%-�)]�\P������c#���ʇ���f7}�t��V/�S�K�P�-��@�S��@D�qT"���w%�V�U<����m�����j�1���
8�7E�^�[ԃ����t#�,&T��W������z��i�k�M�ĸ�������*�a�[��r�����ӲT���<�;�G��o���w����@USq�-Y���Ol�U��IG��m�I�\�A�Vׯ4ۃ��)~D�3��X-����\�Y�2ueh���:P9DB>̔�rVֽ(��PQ�$� �`�,)�u`7BeM�?������do>{�n���,��	�ǭ5����ddSf&��h�Tl�����5/d�>;M-9���i�^��j�a[	�b��V���_����Ȣ��L�S��4�
�,*L2z�)�9�Tt�&C<�#IO���?�ޢ���q�Q��ސ���b:\m�����¸�ƹ�����M�P2?lI� >�f���+u�3��4�?EW�ȸE ����Bc�3+�]&��p'Pմ	���uŴ�E��-��Ы���2^�F������1�S�[R�`�iB�k�W���Ǜ��ŏ�����x���1D=z�v�5lU�ٹ� q����uy��O�
��<�<�l�ч�="�(�e�F��z#ܐ�NK��J�,6+my�zl��C�V����[|`�߽y����)f����[A�*��O���`����U}|䈦�3�m�/�"��(�%�����2���xr���T���Q�|�v��#'�=��i*���pӲ�\ ��8���֎_����#���D�(")N�1�e���.�-Q���l�h�}�H�YʒA�<�%ycC%�B�W9B2I����I��p���īf��b�.uƐn<��(Y�´[Q�Qe�?��V:%(���������c^&Y��2�Ue"Xh1,��􁖏�l��NL�j�Ƙ��o"O�N��79��
���P[=	\�!"�'
�`��eQ���@�����}����5#G�����>@��ѓ���j����jip��ەKl��~�*���47JlM���I}�Ki	k���3d��ILQ`H�Ơ!`Q��y����篌�x4|28}Id�lԥ�h�wi-.�KB�@�:�Z0P�T��GA�l������HF�i�]?�������h����9�Z��	P�g���ԉ֞����Pg=�9�����?�fH��[��tF�~�+�8��hKM��D*E-/��^Ɲr�d+���%~��5&�DʡĂ���\�㡠$��pu�OC�b=����`�������6����.+
ܓ�S��g��&z}O��F�ɰ�F<��:2�~�Bͼ<�����8
�&k��u���L�7iU��e8���gH#�m�������l�5(�w�0�wf���������jY3��L�x��$��`wmҳ�����.{Q�֩�NA:iA?���4a�uQ~�F�l�Ǻ���,��-��6A�x��AJ�髍<��˄_-���V���V��rKY�DD��AT6������%��|=�r;h�m�&l��o ��!'��U��]ɱP��M�fh�#���	�`����J:z?�
V�"�<!_�W��L�q�o�0>������g�E>>K��#��;bE�������p�A+�n����q>��6x�BhR�G�l��a+^d�j0f��0��L_	�v���S �ş���4N&��	(O������1�2Q!��O��.}jV_�g�XYmV�Ȁ��0�m�?�~�sQ����Мy�g�L�ˠ5�>����� WRM��.I崎/*!��ML��^�D�ʺ�{����r����un���~���pi�GO��t@b�Q��l�458�y%U�O@S������X��|j �iU���X^'�\&[�iK�4PT���D3��������7�z��UY�����I�L�S�����L��^����S�W�=�j{mt��=q�i!��~i[�,�C�9	�oN�+��b�P/G�K�6��R�׻U Qm�{i��-h�'��LHa/u�E��Z��0:�L�������K��('�-p�Nq��
���~�qrN�^����N�&��h��� ���Ah��X���������|t莙� %�VnNZ�W�]�w�)�Ӌv���?p��F�t|�T%���Ұ�����IK�]�ΰ�|^hM(����*T�6�&х�=w��A��w)�#�
���5�q��[{��K����[�|�Λ�P_�$p=�ՇF���<��8s^#�2Zr�2
��������G� |�R���F��%����%\�,`�Q<I���o6���ڟr�w�2ܮ���V��o�O�TC(�^v�5�B�Z2h�ݟ�G�p�l�!��DwY�L��4�^Q�^�ށ��G:9����*FA:�s1�''��tc=�н�{ZP���<C,�?J���䏢��UKC��JAL���;	�Qt&s�ُ���jH���O��,���5.������|􋻷�.h�9[	���)��u�L�;d���	�}�S�t9��0jh��Sp�S--�Mq��/���هH��K6[Af�HibZ�J4���E]�ۣaI$ȯ�G�r�(S&~�6\^j�/��$=��Lގ[�[����<�ɌI���y�����XzN��<J�'<�_oV�ͤ�[�J@��>��[?���1.�r��M��ߡS���_yey��ö�=F�ݡc ��T�$f�6n��OSV4R����k�.��wyG74"�P�l� ɻ�;*�U� �}�w���hr�<���a����
�,�������˪�LD	*�m��!D�vx��b��5��X=����eX���~��G9�\$J��I|Pp���ҿ�$���l%-�>I�G��c�i��sc�QY���@cE�;a|6�@���K�]FF��"���B)���2c~k��a
!���mKѨ����w�9��<?�R`�IĲ��D
�ռM������"�(��vd��̉F�2��Cjർ� "� a7�ŏUtx�J��vQ~?~y�������^�Z��Ʋ�]6�7�jV�l�yi���=��,�p�糖sx�ը���A�%ǆ��j \-Bʪ��W�Qg翉�F*y�3�����77�������β{S5I������U���C��t��0��@�u*�z�8n��*��C���� �T��O��.pD~P6��rC�-�b�1�qiYa��i�u�5�^{�c�y�c�C���X@t���7�K/~��3f�������q��]�Kp㱦�(�'ʝm;�/O�x/��sT�o�:���������S�E]XCR�Q¦���?%�*-��9K Ǳ'���0�^�t�ӄԢ��'���'۵6E�g0޸�X�P�kx��JDv���:����6�tR2#Hb\�(p�Z�G��ݓ
�^h�"�sk\Ԣ��>͞����7kK��+��V��0hD�W�,l��%sS���psSf�cg�~�l�琱:؋�j��jyI_�5�Bl+ƭ�d�+�����~Dq��!{Y?���հ�{�<U�_���pA�s�����������6q�N�k�\
/?A���3��nB~�_��X��窆�-H���&#;��ǜM�:�?���)g^��Y`W�>tޫ��*g��:!�7�������2S�G���y~�Ï��Xb_���m5�c�K�*$h3�q�����؟|���<?���!J�$^D�I�8����#W����5{��������QRW��:�b��>y
�P.���2�Y����4o�2d-��͝{�Iy��.�[�k���W����<	)`��@g�g�;s��K�9�jw-y'���*_�G������\C��TTS��Gnu���εw8�y�^��9��6X��l��ov�jI��ZRJ��R�1�RY��K��Eƫ#?��X�u���SX�蓉:~�K��T!������{<���o�@��]�(-���,��0����+���c����a%fp��v���=w?[f��b���׶�m� Wy�á��oq�e��z�H�]J�Ȏ����"7�&����A������$��\j����C\g��$�g���5X���Ï7��b^@D @qsy�O�_#w���F�~�NJ��_����9k�U�s���:���<���ŋ��O���!h�}t:��a�	�;RN���t�(���d�o<�P~��#�Q��g�=(_����iSFV	k�����F�9`��8���v�y��7=�5�?L	Q�����&}��n�֪�$�N�!��ʂ,%�9�>��IF�^>ژ>$�3K�m(Ll�ӖO�! � cf��Ō}�������g&;�?��q���6�t�<��U��s b�����Y]v���0ҋ���:����a��nF�2�@�Kz0� ��@3�x��d䰂9�}N�R��~�2���B��"i�h ��D��1Wj�ّ���mXfM�����.L;f�	�l�����QxJ�^�0�b��@��`�9ZlfL��G__>_��v�^��ƙwu�l��Ufl`�����R
Nq��H�s���4�)��R�#~Kv�����(�v֕�B��Nߚ�)'2�k�2�i���Amփ/��g|M�J�&�+X�����?��!�S�XW��Y�$w�c�n�(��4i���/�ww1iz%�WS8��X�j�T�i����7se�ĸ�vB�*,W�d>�e�A��`OZ=��m_L���E��=����P��<���,��	���t�ù�u{(<�Ɖ��!�j�,���˓�s���}�mC(�NT��ƦP�2��`'�:��Y���#Ž�ǽ&����f��]�(�ji���Ň� o_N*z��y�0g��5��"|��>�8����_�\���0#��r+��:l<*t1�'��dy�ί���B	��� �s��>�S��ɶ�38��!
�{��9��/.�~��h����Á&�F�?�J�8䲭	|�E"1I�e| Jt\`�8�Z�=� T>�'(��Z��#��O��h���u�h�q-�K':.��I��AHP���#�ʳ"�:'��AC�-ЭBxv]�rz��# #�uT���$^�}J>s�}��J�V.kz���z���BW~%s�LW��?����n$��O�0
���l��u��5Þ�d��|����yª�m[άFs��|��kM�@t<�4W���� =C�SG@�.$�0q��Q�C�8���D�����X�O�o'Md���-���n�&G�VW���=+� J�U/.HX^^�SMG%�<B�~,y���]�����46�U��*�~t��3����X�ţ���#�%ԧ�!�ST7��+k�G�5�Es��@7�4*�x05*fƬ]�z���� .��F�V��:���9`��cl1_��l�%&��H��"����.nߒ\�~DHF�_��v9'�y�\���V��,ëC��2���5���ǥcl��8���CB���7!��P�'�����'?���N���)��ה�E���G�
p��]o*����V���~x�������r^�6�J��`;g��錇P�*��N�!p�X��G۟B� �n?�n��U+RC����9�^�����6p�l`��'3�!?&e�>�"U�0+gg�k<]ƴz�{
���Y���uX
��H��Cg�b�)h�h�y�B}�;�����"���Կ�HP���G:Q���b�[��wl���o���?��K��k<0���c�Ϸ�tv����UAJ�Ug�L��/���� Ü����HxwP�c(q�U���gX!��u�����M>Mfx�Uz��P�3�y��������94C}@a%{qX~;0�6�f�)8�h�t�	*o����5L��\�o�Z-��ݔ���E3�H��Y�8�e�Fg�_��߬��r��$�k/p(z˽�k��?�o]�z&�k�sW|ږ��W�-$�O���Ͻ�� >�4��j��ȷ"���^��n�T�ǻy��
��k-�@�^��o>4aS�^�ж+|��/���V{u���p��п}O��٫�z#P��-�kĸ�7pxe��	�t`wp�3�?���3��l���y���Pf��3W�Am�i=���P��R)��Yi ��=t��nܴjT�7��T��Y
~1��/��\+�@D�W�@G���љ��T���X:,��(��O��[h�wS��vSТ���6q��2�� `���PU_�h�LZ��|�E�:�n�ux�W�VL�踀�qsp�@�#�fD�|�Zj烺d��[;y���i�)! �K9�Ӏ:\E�ô�
 	�b��u 
�]��FOh{�P�\�m�W�l(�P�����).�
�b�,ʅ�?�! ���,����Ǘ�VU������*Uh�Ȱ_�XF	��t��#��Fg���H���5J��EfW�ˉ���8�V�Wx�9��N��v�=��L�%g�3t�?�����Ew��՝�D�;$�9��8���*� YgZ\�=l�!�3^�̉Kܬ���&�ExC�%����91�L�^*g�z�f&�%�*�WEh`#�^HKݒ`�*�l2�{Pf:n�Q~���8��yW�����ִ3�Rm)��L�#�(�}��,0�F�u��0D�N�i�����P6i�b�� {^H&W�Iz���]�p��-�k%��`���[P���ˈ4I�V�o�[�9 z|��և�b�傱gs�[ZL���>�W�Hd^).�M��Hj��Կ�cZ*��t����Dx4h#��1���
��.0� ��DG�����cY��V���9r֧��&��$Ĩ!�v)�:\?FK�4"�������.�m���͋��]�^Q�ѥ"�5�FJ;�&�8��Hx�=V���J�2�eD8�.2Wk�O:�:т���xt��B6x��eMm��Ln�	������w�]0TH�^�Ә���59���]���`{��d���E[֋
6$�0�=Ǟ�99����s�X�M4n��o��c���Q@N7��BHn|���j�/�D܄�m�b�H�
E���^�5:>��GlY�c�6�N�J3�Q��8�غ�ͻF����Q����댅5F�.�K�PS�M�*v�m�L-��L�� ���m ���w��;��wm�~@&��+�Z>�
yaBWˍ�b���[``����a��ר�@�y���J0��q�� ��/5m��4�U����ºq�+�$y�1~'=���Mkb��@~(�I�r+�T���G��WD��n����m9��÷ք�\�Y��t��&y����v�pM#¤=����#���|m�
O�y��r��e,���k�
�6��Y͢b-��u)�L+x���~����~�o^���s�����& �=!s� �=�ɼ�L�)v���x5�����2�XEy�tI�������9�\P`��{�����I��^i�.�95�p%5��b@��R?����¡*�$o~x�|s��\{씡�e@�z�.������>��M���,}a���O�\^����'�Y�0;���X ��V��N/Z���g�<m\�z�k 'T���](�^���A�<��;�_������-���w&���q<�M�C�7�5�@����<µ��Ḿ����X-�=������y^C�vʿSJ�!���6W%//[ ��-NB��$5�aty��<�&s>�{�[����ٙw�l4�S`&U�.��)���'�m��y���{�$mr����S	N/��A������SLK���B��B��p@�7��ԫ�\d�������L��4�d����=6�+���|�DF*�[��ظ��3%�H=����S�D�H���{�+�ˌ8�����TӰ�՜�WVl�O�i�e��8�xa�����ዯ�p�B�C5z$��{�N��%�?^;��cl�칆����� ��e  ��t��(�	��i+at;�`�M�da�~F�:g��"R�^��Z^Ǉ"otʤ����\��'9[�F�}|��I:� d�(�#�6�1�?�1��l�p%���T������B�9a~p���ĦZ�=�?���&]ԮJ!\MU�\�Ū ���׬����Xj�@�Ed��MW�����ROB��0��ƞa����e��ؙ��N-�d�E�t��P�lH�_-+ �@`w����4R��('/�U�u��w<���5�b��V]"2hm�ĐEܙ���eT�Cc��e��м��怶�L����z�z�W$[ɪ�����'%�'�Z��Ey�зHIR�'E��%�2gtR�Ux|~MBX���ƙ�9���ߝ�FR�ܠѥ��܉��J1$�����*��
]��*f�	���z�Dqn.��޶��Jfږ7�w�� >����\���%���M!��M�%��ז�ƿFUj���l�V�~#�Ibv��"�TF)�b,6��c6����y3�h�d�Q��ݒ��`�@��;��oZo�R�e>���*σ�.�	��Ua�����L�V��&������,�{���LSn�b6pHa�OcS���C?8(1ܥ�M���=�:�c\%lQ���h5������ ʅ%�#U��O��{���D�͢~����M���5dVۘ����/�D7��~�K)����d��h٘�B8AI�=lK&���7܎�,������Nw	�eSĉ }�E'�Ђ �=��:..o���J!�R�o�	�~�.��Ofo �:>��	���0�+�9��Wtd&�J��}����������tɠ�k�-�~��xy��ڄx��7y���]졈�����h��j�Ɇk���5�qI�K|ǰ���NqԻ+��B�{�)�GS��PpB�y�!��|+�^�"��HQ1{���Pϳ;�R�D5�?�N���g�	�	��ݭ��^�.�Cر�SŨH�H��/�80 9��u:�������f-��
lB����¬��-��&�����&�}�c��B��4Ol�:윕7J�}��t ���r-����+�`b�l�1S��׳ѡبҟ�!l�i�G�Bd�[�^�H��D��6�$]n]PJ��|{l����􂰀���3��v ��+|A߲
��d�Ir��z�jwú
y���uJ�	�Z�(){���Qe�MGXD���w͟������:e�P
��ߩ�& �������+�Q�%Ǟ�(0��W��UZ�_'�w+�lϼ;x�/lBY�>̼�=�h}����n��������$�V��kl����4�,�d'�g��.�}�:�,���N�1�򈧭���1>�-��<��M�G�X��C�@z���Rv�Z�U.�Q�MĿ��B���<Kdf������+8:���m��_���ڦ��V��@�4��(��xًp����iY�����D�Z6��G�zS�|�զ�>�������E9�]�W��-dR��V��>K	 �6�%��M� ��l�,�/��KL`>�8R�1Cn������T����E��!��F�Au�����k���)&٬՞���l[X$���l������� �!�#���@�7:l����jO��ƇPx�}��ƚ���߱�˿��}L*�qEX�\�Tf��e��N3}8����(<.:Pd��	�˯K)Kf1�j�N�ŀ�ꂣ,.��
8Q�׷�ן�:��>�#i���~{ؾ`��ޝ�J�q�i�#;a�g=W(�;�5�T-���
��?�4�S�Vnw�^������?ڃi��u��h�?>^������'�W�΄T��۝'���`L���{-
H���h[.Ł(<�t(0��@r�|{�eG���Y��q�N�f�=��X׌v$�����+5#sԊ��y�EZw�_GQX,���{�$H�+a�_�GO�#�v��!K{#\Y��w�jb��eǷ�A��vg( ��:��޷�Y�� j�ev�uS]�.Vi�drxz�f-�Ցd$�A`ɡ�
s� �����\��d��W���>���T��;\g�&�|ڲv����(F��1߂�1�eB/=t�5����d=�y���b;�v��G�"W�ҿ � 4�5D���/�B��ú��e�$���ź���)�/>��ۅf�ثx��_ɾt���o>d�f�r8�b^��f����\ٙ�L�r�B�^O�֞W�疗jH��S<5Sj��1ǐ�2�D��K�=;B����A���r�c51z�������a��p�dr��X�$��o����%}���F����Ab�R�da>C]��P�%�ݜ�@��o�A�^/���?��`nh�C�dE7�Ux�J���NP��Sɘΰ�5�Uqx���3կ�xd�y�P�)�����Nr�Zj�$�`pmz�0=z�,�6�O�kp� ՗St
�X)@u��7����2ey����@Kr>��O��A;���=�N
p&� ���M��_qwK��V�؉;�)� (mF:_�Z���|iq�oQ�\3��2�*:[��yș�Do]���BtNDz¨Or������f���؏�CK��+tC*�&�t�y�"q_8�b�|f�������b���J�Hn�i��SJ���Q��$�U'٧�k�"��k�)!�H�e}:zj(�c]�>�{9��ܨ�D��
� m�*qE:�;��f�l�붿4p�!֟�ǫ���!����Z37�����d��½�=��Ul�8�/�u��UD4�i!(�ـLrL���V4�C�,�al
�_0�P��r��ַ�����B�c>���u����#t?A�$�o�J�gY�pP%;��k���f/AmiU�|8>l]�ϘG��+t�,���T���e��������xX.�0����z�~oU�=,Ɩ-=�ן�;�^q����
�{��bҖ��I5Cu�a�Ù�b͝��>QW�;[U�-/��.S�A����<DJz"d	�>��ZWI(an����+sLӀ�4+�R�I-�ٱ.��H:���L�:~���->C�>�lb��' \��8�"ʘx'Y��R���~��mv��c�UO_�<�����^쇪��s�1Ds\4��p8D�]N��A��R�~�|'����*%EK�dJ�f2S��kXY
��4ư����3�����y�������|y�v�tq�,&	ٯT7g�3�ۓ� �@Ϫ�����>�ߴN�J,{���c�������W8���3h�ՠ\�u;PEnv�^r�>� yA����Ưk���חꞒ(hO��˽�[���b�
�b^�����p.#k������w��iyDBG��������$�˔IW��^ٞ�Ab^>�m՞�1�R�!�	�#���ɽ�gC�:�Ň����a�E:� �X� �az�Q�UeHۂ�OC�8_�o}>]�x�����?���t���kxJw����Ǳ U�� ;�E����;$X��B�}�u����Rn�v�v1�[��?C=$��əC�=h�^&;�=�T��5Sn��ɖ�@J�����V����\�gt��;3��6r��\, c��xd�]�t���rpa�B��c���F@�y#�xo�D�=}r��>.-ӯ�emǇC�!�s'/^o-��+�TEXN�����A���!�U������Ǟ�uȑ�A",�r�E����&QW˽����シ\y{_I�IW1�:	㣦���Gv��S�"�����,#`O��nc>��ݯ�q�{�Dz
`ٺ�>��ߕ��k�e<vX�o6��v�όgv��:JM3a��l����S�G�#֋��{�>�.�F��KbdteĚlջ�^=x@�&}BsmpvC��	H�� ���Ĕy �F�JN�;�j}3������{7]��S���p��Y��X�R��Pη�<�5��7s<r$`��Z��#��a����ǰ9�R={ѳ�5�f�8�]����z��R>�kT�;��$���9��H����O(f�:s���ul����XU�0-�#P��m��cY&w_o@�'�Kn�bfg&�52�D����K�!��N��!���l�k�x-E��<C�`"/z\�	�j?
��ͦ?]Z��S=�����aǳ�SO�*�E7�u~�'zLn����ƿ04/-����`~� L�׿�6\�@W���^i�έ���w�łocz�N�d��S2�"����I��WyX=�=JhJg��'n�9�S�MԆ\c��\4��׋�,�U�c�ωC�t;\�>f"4u�9;�~+���a�Ȫ=(�	~��������a�by�m��Gdy�����ǵ�&����/�X24�F�4}l�,��	�!WӤ���h���h�Pzr�yЍ�G,��&0�$6y�j�̟�mk�(��4�� .[-�>�ԣ�_O��۪n��"�Nߺi�9f[��)�G~��
����(�Z��E5�i�T�U��lࠎe��[(K��'?Kh�������;n}?7���QJd@�S^U����
S��a�֠B_�Io��o�<��a�B��>G�L�G�By�������`;�o2�F~Ҫ~���H��2�m��-�z��'���H�(�&H�BD����P�Y�����|��A"�S���Nڳ�������\���v���a��KD��S�l����fu��S..CC�k��0�S�*P�=]{��.^��ӛ��;�q��h�͊���
`�� �<�2kq��P�)p�q�&��m��ㄜ7�<��%�-�%󆭼��2�������6v���綕�zi"ɭ�Mu<���1�O�;���aRj>}�.K��jb���
11w�_�g��otpH���V�8�X�T�5��u-dZ<*5R���2y[5N"���O��:� ;�y�a}���!'
���Ay^�&܄�@�w8�5�V=M�+�Ě��G�����G��]:#��a���%0����M3�;�yk��k�G�R�}��c�y}18�,�p�)����ݧu,�<��_C"��qR�x�dy�D��1b��a�o0ԭr���5� ���h�.!zjGC)�58���Ea������~H&j�z;`w���X?}0>*���6�(3:u{5y͐��U��9p5�T�Q@�3L���<č����3�/��C���1��nn�y�63沠
�����8k���?B���)ؿ.��O�?9O��2Y0Ś?�Dְ���K��䉬p#��_�b���Wq@�Ap�Od\4<��#g����Kg `��8gkei�u���QVXm���/I���+#o�����á�rF ��P)�m�ﳞH�{8$#�Kj�5��D�JQN���9�����1C'6�f]�d�Q�4b.dl4;���4�t7vk[�w�Dz�t�����T�ز^�L1�e��fܶ}{qB�������%8�}�y�
��wC� z�A���
L��p�R�bd(��o�YI�:�03�+;y~��7F><�z��^M�&M�˦�ٴ������_'ݙ�&ό���>6��2��0c�\�j�������s?��R3��Vц<� kd�g��M����4��R��We8��Su�C]��g���Q
�"Ep#q����n�2,�8cOu�Kۺ�����;�L`�P�{E_$=ê�j��PAE4�O6a�Ҍ��"��N�a,)r�7���rǉ-�h��XI��˒3��]��E���^��@��j�oap�}K1 ���R���S¿u�9�� S�'j����o������F1��(�zM^P�����v�s ��W��#%)O��0��K����0�}��P��7��{���*�ȴ
�|뭲C�u�خǩD?i��G��~��n�{���T�������V�x]׍�7+a�ä|T��.mC"{i;�wA��n��+H ��Yw븱�*�W|Yi���%2��|.��T?#��"���[j>5$� 6rzp�'�m{FM�/uv9l�L�
��X�m�\W�%�B�]�RZ��A~V�{4h}�,QO����J6��,_�29���6�=��_kWDЭ�t��X	ph&<�s�r辒�r�k�ީCa��T�D����;^�Oj�� V�2�S#�`�MY%K�ɊDܙ����P�%�Q��d�H��-"!���u�5�#nv����Kzkx�C���	���V]��"3��y�nT��ֲ���A��;7	�����(|/Ͻ?,��
����0O(�D��u�f���|�r�S�Gz{.'d����c��;�6fX���MV}�c�TZ��[O)J)���õ��:׌��E�9}s���\	�_%��#AԘ��8�L1��6�]cFS��z�ul��z�5쩏	n�X�,ɜA;0�W��z��fu��xh���*^V*8-D�u7��h�U k�ڝ&�� "��vO�0E6���JS���$�)�9�ed�I���/��xO`s�D����)�!�d�$��&�$�ˬI6z�a�/�RB���F�MI<ҙ'_#Մ!��*橨���Å���G�պ"
 %kJ�ge&���������(�B�x�0[�/�B,��� ����X��,�Ce�����R`*�i� /�����Q=�>�����ܿ�����������]<��ۻь�F2��(��T�g�!9IV��o[�RZ���<7I�)���~�� �0��Ad*�lg��r�e����_�f�h���r��Br���c��+J�<��e_Ȓ�d��ǂt���?k/GQH^=���Y�h�L|l(����u��P�)�%�w��S�@`�� ��V����"I73@�l�K�ў��5t:)��'�Ds�\�.�S�I�s����#�A�O�go�w�{���<�c65�Ѡ�Y^P��t&z&��Gm3�n��\�D°��ݝ���$Hؿb/dA�nM#������Lu3��1�롿a�D�tK����z�q�/��֢�ͩ}@>��)�Cb�2R�����Pq�ٶ�
J�ď���l�t���\��D�<�[���×�0�!��$m(�)mT�].��,2�"[�p� s�1�*#0F�8`}�L_��&������]�X�m�p��b�!C���@pnP�W)�F�'f���T�?L��o�zd�p3��3����b�$]�sC"*�!���U%�7�CS�uQ��+�@?���,��O�=`�Cƚu��JH��4�)����[�c�	͝E�"�U��u:D08E���V&��3s�#�� �fNM'�؊H�=�����~ی�~���8��j�>��� �W�n���v�QH!�f=,��3�g��pn������ !Si��g���vhT��`�o�;L<�9���"@�	.ȷpMDJ�3t�_��/Ŭ_����`_�*(�c��!�O879�:Z`܉1�_'��NV���oBX����OP�I�ǔaN+ϝu��b�����C��,����x���2�T���jE�E��[�g_�o�ٳ~W�Hǩe�D�Gv�1�]���c��[:[F%4����S�*�]%���b̄c��7��ߣ� �}Dǘocߗ3.h�ݤ]�m	��2��x��t�@��4����cs�{��St"�f���)D\�ΐô�,�|��L;��e���N����i,�UԘ�"V����>l�Иd���p�%FV'�6��4"�,��c C��)�@v�>�m�ջ\~Ӳ��q�9��܅m��):T�o9�
���*�fɄ�6p�E_ǻ�}A��a��<���d���D���Ԝ|�`��=8�1Ma:�e���sx�H~�)�ĳ�V��$w>'<�%p�����<l�x\JWZ���B����ҍ�7�U�F��(��-2Ͷu������� F�'��1������݃���5\�Z��^�F	n���ŗc�Z�ݝ��x"�*S\pZ��.�p�W�섥�Gȡ���|#�`X��ࠚ�Rs�C��SCI<��C�X���.X��88�o��Z�p� �qݏ-��yظ�DEH WeP�=i᠓�"�ߠ�r��l�ɖ����_C�E8�����ZLA�X���eq�\D���i��/|խ2�����(�������x�5��D�<{r�0�UM�ѿU�H��w�p@�����y}�]G.�%��	M��O�ܱ	w�A1�[�凜���>��J-<����8��9Vf&���]�1�ϵ�D
Ȗ �
��� a]�a"�5�U���C�hz7��-������s(��|�I^'��d��t�-��`.ƚr���EG�"��h�n�U!��Z	@��]��U��U�Ԅ&�>3�IT�1�/������,15���C�h_��p�,e��W��Bs�k* ���"��` u�tf�ȡNhLi��W8E�
�Rj�n���2�D^�N�|�W��{���1�3Af����ۥ�#�+��$�8 ��I��XQL��Q�4�@�����VS�A߄Ǣ;i\Fi�-��f:7O��j*�밻s�� ��k9h��8��xC��C�va�,�\��i�2TH>�0���9�c�#7�g��s�N�T��%�iP���Z���M��a�����^��������IQq���2a��6l�^��3Ƀ(�VM�gz����/��$)p�9P?*V�=p�fv����:د9'�:$���U��z�R�7�BH�ƪl�/U��fN��4.W�2`�����q=|�e]�%���$槡��a����1R��.R.��I5(�
�@p����e��v���9���F����_�{(3�t�Z���TG���=�C����qwHL�*�M���Ns��ֽ��;�����j[tF�X�c�C�XL��'�����~@��]sPmO0g��D����wN�ݕ��-/��γ��DbXj�4X�<��bh��+�Z6�g���ä����L�H�U�9��Q%��즔_�w%�QOt8��<������E��|�\h� �'H�|E k���������!�b���c���?�B�P�[M��~2G�G�`��������7��u����)��r�B������&� yO��e;��)4�Y�6^�|�o��1:�W�h�g{���۰����Џ��d(��%�1�ֻR�W%�@J�0���YQ ������������$�Lf�I6��6<�jE;��M�Y���A,"-�"�p�w��. ����3���eS�T���Vi��.x�t2����L(^���Z;����e�x�+$	E��/�C�"L3P�dڌ*������������+ �,�N�;͉�t|-�sj�[�����/��S�` ;E���'i&�p�58iUH(I�뛬���U��'�]j��+��T8�V��hJn�ˆ�����!Mn���[C�;�e�}$}����2q���yO?<�s�qۨ�//��'��5D�w�1�o�Ϋ6f��ڋ�Ǟ�g<"��=�bd��h�=a�Ԧ0��.�M��RpD �&��m"�m,�D	UD���eXo۽�+�$z7r���6����U��K�e��'�2dȐ���qb�B�!�bko��"o7܄ﷄ�S#���ةJG�fI�w�ڣ�C1�?a��B? D���cb#YZ ���OX����H���b=`���F��5�?�^ s4h��		���e�-]!����J�]9R�A4��S�y��5������z���<Y�7��}��B.��]��L��F"�B�[k���Ah�;"�F���K#�Y��5F8�Ia�M�#�6����'�^�/:�Q��p�'�-��Cj
�  ��T]H��s'�)^FZzFc���Ω�.�H��w�J��d	��ls�۱ �s�x{k+\y��%�o�}/@΍��m���u{�c�	�i���.��D�B�E��u�����F�j��[g.�{��Ug(}�u>�ؼ/������S�w���f4=�}���9���s
5Uר�b����/��*!-��W�BpI������o�#�O�n���B���8��<mJ�^w{�lWz�^�I�'fǯ��>�-M�V�"Bxf�H�|��搸k��s���I�3z���W�~���	�6^�rR���Nͺ�i��&�r�	
;9U����D��"9��WX~:����P��ʢ�t���#����
c���0�a%��ĥ�j	L��Mu��su��gFsV9�!휫\}�V&�{�)� ��.�t��߉U��G��r�Fo�jn=h)�<�u������Ө�ψ�A��Xݥ��l]�+�	. ��� �a���k�D"�'�T��O���6��?=b;p��X��b�<'����/��L.�,�E��{�8xx��G����!#1��"��0kk�Ņ6Kn�F��N(4��ZY3j�"�����H�@`[�[��.Z�5*c���{��>]�iDIY{{2�G%-�|����A�N��{+!��"tL�$�ă��;*Fw��u��1=�(���68;3���{�����DLY�%�����-͟�u�R����4��p4��ɕ��r[�l�� �4[z�=Ʒ�����t�����J�3�onn�mC�;�yS���U�r;iP
�*i߁�4Z�!�I�7Û~�p�����e垮��nA{K<�8tL^���և�����5�O�4��=LaV�ٝ/�rY��	=�xK�UTb]�ۃ��o��:����Z�� V����~K�0u�����'��Q^ǟc��K6��q1�󪉎P�i
�΃M�008�T?1*Й6���h�����ۄ�_.�Jc>�#2��	�̜��j�:��ɜl]Jz�\���nZA�fp��P7	�0��c��5Gi�ܚ�^K��o�.���.�,06�'��N�.T.���y8������7����!�7,O8z�p����~H��%���9�D-��'z�͕��
�Q�ePf�/���-����������<Uw��E,�Tr5�A~3Jf��L�L���,��t꧎Ӑ�����V�`��2�Vݩ�u�
�ݓ!�s���P}�{vݱ�~{b)��eG	�-+��dCR��"��Y�������jÇ?w�K�!���zf���B�-���4�m�~��_ۇ��U��Y!�:ܭ�+(1� 3��ĎW�m�'P8����S`�-;���za��>�H���ծa�$���w����h�>�[c.zR�fy�ō��w�r��o<�� ��&�Q���d��Έ! M��8=8	�t����k5��>��Ӗ ��H�|�n��Ȱ�]�a=�)?9��Ě1�ø5ph���~F��J^��Q��P�Z���4�����ǝ�~I��@4�l�N|��G�< 	��UoFт(��r�Z]Ȩ�^���6&'�ƑL	�Q%�&E�v!w�W�� 	Rt��~V�"�]�~CՇ����FuJX#�[��-9D����5D#5�z���_�8i�KRA	���qe���I�K�i6�U�ƴeb�����:�s�b�`�C��ΫcȖA
j3]�|�I����=�D˨���\*�8�� �u��ҭ���w�ړ~�������ONF�]���uO��ȮB�+MPx�fc�7_����4�u�o�?֦4X�YӼ��r�/!B?^}T�����������L�ڼC����3�����Ҕ�P*[Ō���hk��H��:]��
�H����Ѡ;; ���d�ԓDw)�������F7��ڪ�B�h[�L t:"=��Ӄ�9O�Q�Z��r�I��Ǔ��F���SgX�L#��`�x�S��flU�%uۭp�l����}M[�/jNX�#�!���@,�:Η^��'��FFc'Gx<��їz[�O�� �o�|W�/I�tؾ@�]��;���7ӝ��AR"%$�~98�+%�N�S58�5&������Kꍅ��0���Qz^�>��D2ķcq����B�Z�>q��S�_6�{ZW��/���ǁf^��~�+�8r�'��,;C+;.vl�n@�Wm<~}BW��#�S�i��I���_ƌ�*XV�����J,
۠H�|�2��j5�a�&�}x֥��X��Q !:���(+�{��N��x�z���*��i����}���"��P�����$^�i<Hx��$�o�ҍ�c�ya�'�=u�C�*2�dC���j(�m<�u�Z�=�ӆ��}ߘ�qQdw�ef7F�ae�'w�AL!�x��n�!�(���5����t�܅�V<U��R�� eb?�[��0	����)Ha�s��ج`b;��z��ٲ�G��\����꽎3`/�.79�^�(L��2E�df����čo>4��¿t��B��2b_�gnܪy/���[Z�&*B==e
q�H�6C�uz|#ć?�xz����ƅ���8'^�V{�n���#��9B-�J�Ett�haS��w ��Sb˵�9cKe�cg2]1�\�>Q�~�z���4zժ�;'֫�	�C)cCn\%�b�ǽV��3���zԾkYƻ|�~���T���9�|�
�۞��l�ڎp	帋�獺��q'+�:c�J���	�H%��]p$F�@�@uɵ��_J������q�*�⮀~�	egx!�-g�c���v�;�#�h�C�� �P՜�Q�<�W{�uKQ��nv�_�퍪%ѯ��0
�#I�J-�ޜ���?�{���h����6Q�,��G���ץP�r�!�L[����L�/.z�U�T�Q�m|ϒ���R�c��*_�A�����k����_�PAh�O�4a䧪��ag���1��c��_f�k��=S�]��_�n�T1](	�j��跲C��)M��@J�S�����#a\l��+�UQ�U�ý!��J!�*>2����/��"�n�b��v'q~���9�&g>���{�M��d$��c�sҨuȖ��.���\k��&��,Ku���}���A�pՕmJK�%}kY��z<��L~�T�:� -�\��,�������f��	[\@�9f�����d�h�,,�=��ӹ>v��E�X���>����g��h\Q�]�؄��V�}N�>�QR���WYu�Nӹc��]w�X�]<u�9wa�rߪݱ;_��!��Xo�8ߖs���J�!O��ds|������[r��՘���Sz�^囈(��.{X���U����|�G1t#�RTosq���8S�٫�צ��٩��r��3�Aћ��V�0��;�a�!�>�,��\f�)
��������& �7ώ����p��sQ�:K)�"u�/&�>���m`�"�Y�bz?N ��е�2���\E
#G���I�7�������E��S��a���e�$��_�Ŵb�]��.�v����U*wC�ͯ�^�Z��ݥ�����,���1X�4Ț.�I�~��ur�7g[Um��Bw�`x�X<���)����0�w�Y�h����(Bq�@�]��3�$�!�
�JfV��#��Ų'�	�U����\�����_���V�=lm�&ķ*��O���C����;t���l��U9�q���P�Ṹ�QX�� ���d��ޮ�MG�D
����[b�B#L*�]��X��~���Cu�C��j�<8��F�|x�X�+��Vu+���7�]o/�qE���N����q�C}��o��#y�=X��S@�LT�g�9��4�H5�,|N�a� ���5��!�k��7?ɢ�?�Kl�����Dr�A��*��qH,D�o�7�La�ߋ�����>�O���T�#b��d��~-�����0��t�W� ��|T�cj�_ﱑ.3�rzV9U�r�������݇�i��|gR+�K�=�N�ې�x]!��T�A��N*�.ꁢ\
?��G�y��7���pЪ���0�>Fb=�VP�n!J��V�f<����,>��"�?����?]s�;
'��~�������Z����-#*#��eRF;�!�^`[�u(G���YQXQ�d��1�M���2��t���c!��"���0�M`�=d�ܰO�/ȅ�co`p�v�L�jʛ��U8�Lp>�4����n�[�+sg��m��X��%���]LC��0�f��1����q�Xq������w@�)	1]���d�{_�ʗ��OR#�B"Y�
��d͸2x������:���M#y5#�թ0Ax2�F�q.B��������7�O\�*�2]3�^��0ڼKɰ����!�)|�OO1�����Xر��s�>r��� �������n�lM��:���q��i�!�t��r����B�&��gnOr����9�vC�]C?5���t��DeJf�D��~�9��؈ʐ���
�['p��	2�1�u'���g�������}C߮�=�wJ$�-K`�Z��W}�����E8��xulq��jT+m3?x6�����IB�@����9�T7cuK>�H�	�5Kj�*������P�r�c��ARF�@S�j=�9��F��h����d�\8�8d�#��-!���*��w�U�>�Z�_�
�E�9�~!JJ�����]�WfV]>�lr�@��'?����ќ���$�8:M�b��P�X�n	��\� �wdVug(Q�y'&;ی�pH�>���d`��	����Z!�1<�pYѽh
KEO�\�D`v�;�5�]c���+��M��|�?�����$Eh0����1e�$�sf�C�0]�%p�%	�c�6,���Z9���\۱#�ɍ|4�����IS~F�[M�҈�hr��ˁ��M]�Rα^�E<�y���V�@�ݩZ_[Π�'��{�-e�E=���g���k�>�����I�i��x��U�Cѕ��x�E_�Ş4��f�ռ2��]�ۇ��i�6{̦���f�>[��٠`�6��"%�.ŏ���$Bc�E[�6�	���D�������7RG�~
H�yIZ�'	L��y�pQ�X���A���ꂝ�m:��7�hdxn��A�E�������/��Z�y��RՑ_���7O��INKw�4n��N�0e�7��e@D���&��7���&���Z�2�,M������zv��O�3�]���+�ɣ��]��HM�T@���i�k 86Œ`�PU�Lϻ��nc�j����9�����h�(���?���	�3�>�M�U��|��H���蘚{%�$]G��Y����3���!qL�eZޑ���ڜ��,���AYWX���TtK"����]9����E�C4��B:��
ɗ6����ξ1#3��o�}b4��n�������*��ۿJ`��j{���Mڴ���w
|k	p�f�⟹���%sa���X�D��ǔe�dS���:�a������N���P�E��V�Q H^Nb�}K������0K/3�XR����x��ksO��s'X)���և���#��m�B���"9�e�~�i��p�1ͺ-s3D�P/��L4�.�!�禍�)T\44����thMk�j�b c�S��B:��c�<��v�!팟�xSke��c�0n��Veo�����/_��9��1v.q-��Dʮ]�=P��#$($&�p��3�2%
��z�ĕP����$�%<�S>5�oY8K�����nV��b���96� �0<�����φӈ/�8��l��J�}��2�Ake͙�6�[D���M������_�ڡ�g���fq��4�b��I�!ɀ3���\ 5�C������n�㙾�l휔�㷻��;���{��}5?R��(f��a ��;�#���;�0GN)pwva8��(� �B���R+i进OE�w㱼5\��	6�eV8�g
�
l���O�� ��٘�X���9WeRܨ'͙p�>c����m��&H/�������|+��7n&������tR����O�o������K�5OmE1�|�D4��|���\�POާ%He���6͟M�?���Q+fr�IӲ�g_N��_#y!ā2�D�`�}l^�#���! H`���S/9_,h���m���`�7g�S2\!��+T���5y�m!����0=�����:��l���*Ⱥ��t��3��[Ax
�U�lWi�t��MТEr�2a�Y�<t�B6a2�n��,xYZ�~>)�ϤY:Dx1�9�P����@�Z���t'0c�"��`�՜{q�����T�Y���x�:yH�!3H�rj���w�KN�c/��2��Ď�W��8e���K���Q0i�����莤~s���
�e�6�1�Ra"����..V1�˹�_�\WI�,QI�[��}��) F+��O�9K�.����#���	�.61��h�H)�d�|r�O=�x(��0���C�Ẋ#�q�7`N[�ᮞY���v�y�����K�%Q|���/��ggD}���E���ݝϑ�ވ	���|�Vm�Bͮq��߻C.�mSz�xZ3���i�k2k�$�,��JF�x����=��*~���v3����5�*o���8��Q�ڎ��7[
Z����;����A�?1�~��G�܊f�!��z�qK��GTG����b�]��o䏗�J���K���}B�N�'ktȄ-�GO���!u>��7Ȟ�6�qi�j���o����ܠ̉%0ְ����U��\�E�N@S,Uh��~��d<�  ��������Hn�Jϙ���u04/�Dw<Y�ӛQlw/(���o���~�
q o����%��)pw�b�E��//��e��zxN���T��Nߊ�����P��AS�7���u=ʲ�@���KB�Y�����t"^��0�u��>\k�J���bxY��$8�o���og��!�Xcy%e�٢�v����/zU5�����'_���>d�y_|vR�DPV�K~��t�ڛ��v7Įǈ\�k`��F���e/���<�ⶕ��Fg���
A^O&�q'�9����N�C����=c`ۍ�fµ�w�*(�Ro�a/��rʹ�|�J��r��GMMg1n~���Z��6�sˑR?_�rBUR��p}�e�g;P���~��o��eܧb"���G��p�N[�����!3n6e��gGRI�I���sڄ�0�S����0��[����Hߴ��T���+/Э�f��䶂�ߕ�����\WHgl��ɤ��H�+wJ>�@��b�CTo!@���JL�/�I8���&i�Ď��˅���vǟ�-i�r��q�i/tC|�Ǆ؉�����!�r&�$;��j�f��p���у�+/^l=�\�~&�1I�_��n�V�Ԟ����E4t-GOJ�f�-��ؼܫ|k����mL��}Y	ۘ�u�G'b"�؉W����g2�4�i�,Z��Q��k_^�n�I�S���Fk��w�ߓeD������ym�,�è�fZ�q�5f��%��#|���/�2Fe>I#�y"dP:��~ގg�V:����&�ce�]�+b4��T�^��l�ܓ��Mql�la/y�o��q�{n�7s��׮������q�h�x�����$����G=w�b�ൎ�K�\\(~���69ir�0ew�(��6�)g�]v�ah�>#�OB�)�����.��U2�Q訩f����Gߺ���G�综D+-C��ԙs�0:_X��a�I�H��<e���L���`q�/2CD9z̦M~Q�ܧ��]>�
*(r?Cq����۸UR��v�����
�� ��1���\ �%eU� ��h���;���u���4g���ԁ�?��fN�	<C@�m�-7N�:��oq����̓� �o\	\
���▋����<7����H��^[�t&|<L� ���NPƛ�yqt~Z���:�@���=��Ѽ���u!p��`���1>Q�y|��Y��C����]mbK�d��7�ǖ/����H{ %er;P����O`����{��p��^yփ�,���9y ���`(<vt��s��J����Y4�&&^"�,n�� �����qI�T��2�+�)�0���p��MV�*�w�e|��G?-���?a1������~�9���O�[WSڼ��X�1������ҧ������ Z�[i�:E����JN{	�>��Zn�p�LW�>[5o���y����"�}	u�p?�P�e��X�y�� n�0�����7�\4��V��wn���j�C�:	T3$23w��Q^�ُW���ӄz@��^�qv������dq�.��p���U���-�>�{D)��;wNl�3 !Y@��vyخ�J����ݯ�g��<�u�g9��nHn����
OT���/��rt�j��O�Zက����.��&˝C���ä=���K�\����7���mk�.D�(��(�Ӟ}EdQx��b�i���m�3 ������bJ���۶�	y
�ݪB�\yz|��YǏ�!�?{��;�t:��p!]ֹ���?D������f5�b�3W��zt��`�ЛX$T\n���؆�L�<k��w<�b����/E�����M��cC^"�_w�CJy&�p�STMT��u��:��l��{��2��7��1�����=-�Y[z����6:�v�D`�$��!�s4j�Sz8���� Ϯ֝R""��4���1�W����j��MF X��� ���)'�U��poN w�x��o��}i�Kn V�kz8�f�܈8�&�U�P�w.��@aI6�$Z�$�V�c�J� /S]T�9!�?^3b�p���q�ѡ�yU�n)�s��c/�DXY�9�oԆ�Mc�f�[,��-^k $/���\�]�*���`w�;����9�</��횤!�`17�B,OR����wA�F$�]���f�`�gΤ���WS�����ۄ�fW��s��Z="���VA��l�T������A`�?��{�����%�9���_s�#c���%���Aw2�}�7���  �,/����j�o�-A��ra��ڌ2L�u�-��箾c�N	��'�q�*ʖ���@խ9$�%�q��o���X��5��G?P�i�i��+>��=��Z�B�4ʠ�ķ��ie����]��<𵴖���B.+�ё���~U5mT!]��3k��h!3G�C[�U���Κw%��[#��2��sY.�%�aN����@!��� ʤ�%<	�R��H�I�q�j��0�@۴@@�s�2�;K���E05�����dγQܥP�z(�n��Œ��f�*��G�s����t@"p�9�t#��J(��g��zbR��*0P n��+ ��tqwc�o^��U���+�g�C���Pqx �9�*�����̤�YeY��% ���2���q�(r��?�հ����u%�vз��Ǳ�;�ʝ
`b���@��
�����q�|���aZ�.���;�ŵ����톽x��CN(���pk)蚍�p�^���<b}�S���A��`�0����g�����h[��@�\Gb�
.+n�*
�$3v�#�*��lߑ����yD�jr� ]'�\*PW}�sJ~�;ǳh�nLF�m�Mܟ�k}���f
]�h���ai�`�ә��"��={�"�n�*{sb�{x��HwW�6�!&�l��@#�x�Н$�U�A��v��צ۲��:������.�Z�܊���7^�8Uq6�o)�OA���	#���d,?:py]��7���p`�%�/������&O���l��qD\�e�
���5b���&��0��H���xІ��8��P�3�#k�#4^"�eE����(��5��|���+1b*j�� MX�B�)βѤ���$�If/���
��<fq;"��(�5<�)���Ϝ�^�n���p�ɫ�g5��]N8}0|c u����KT�I�]�t
�}[�:��e��xV���1,
���k���uaO����%v*�%=լ6ʿ3(f�l���p���%��c��a�aE�T
�w��s�[����#�������6-�����x��㇔�3-���@��VL��2�6]�V�li������}��{�@Ρ$��D�ۯ.D�l����L_]O������+}7�U餗���`���kӬ����Kd������"��z�^S�n;`����C;1����9��P�x�`���9�>��)ל4�}��:��PЯ�Ŕ��y"+㏯�D^&c��k߰��x��_���s~�׶��;�I�����k�������uBD��^���&,�tv/S��ۑK�6��>�~����B��4$r	���V�q촫�8�P���K���P��J&Jb�v�!��3�U�1�'�;D�*�)��H��
�$��~�^���*��2�E��ٵ_��,����#UT�Xȫ�%�O��b�P��:�ui��\]���)�Z����t^�ĎVQd٬9γ%h��q?���૆^i�ʶ#�}���V�F-Y����ˋ	+�ww��u�Kz��0h�pl�6>T7�Lg����+$.�����8� �p��lL������ �#�C�����6D�E޸�]��N�Z��*��B��'�N:���p�>�+;��-]�8�7]}\��W��<�����W1Y�q���b���a���:"nh�0{�?�9C!OsE)�8����9L4�����������$cA7��w�[͸���G0`�vp+�Y�w��!�=�c���Ԟ��:ϋĊq�+/�^]�Bs?��7|��JnDjҸ.�y攀,�E�^�����
U�k� �(�U�X�{]��E�^���:��a��9Y����$�,�b������L=��J�֊V��7a���-[�~�q+�R��N�=:�7?v�㔤�'ڴ�l"�z'�}����v���qWn	)��s]*��52��I�At���e�n\�gꆍeS���ꗗ���Ro=�]s�2�ա}Q�J|p]���.�d���{&c^YGԡ읡�>k���H�Kw��<N�m�ׄ�(y��psR�2�k49���[����m8i'N���n����mEԲ����>ӃI_�Ɣ,wNX$�Z*bOav��/��w��/�G�mUv~vQ�l����v��*����a/i9Z��EXv	ϧi��gƫ�n^+~��e$57P@��d���'��A�d�-�E������#�ܗD�sC�{��HP�e'//�����F��%�^L��1���K���;ˇMe�p�}����]��ڣ6�J����`o��U�S�U�AT��7��@_�db��k&�� �J�pP�s���s���1����(~[)s�II5pS�R��V��"����@�R��Z�U_Ҧ��l��F�%&kr��P�X���~PU��9b���.��ޚ�Ml�!Y�N��rj�gh��귡*my��m��̾椕���%,�(�^��~�6�l�z_�0��7��ݟ���>9[����+�Ju�_I�qN�"�01	�n�_!��{��P��Qm��S#aw�c�X�������0��zl���^�cg-�w��&&��)5�4>�pi��*`�|!��ER��Q�6��fIT�v�6�B_�B)�as�����~y�)��u� �"����vA��Ѭ+��(�ں���˵���%�G��	q��ruj����i�m}��T/�R;�*gћ|"�������O���.��zuAqzu�?�X'�+�)�9+��vp��l)�?E���ĥ�����9Q��4�.$�g���rۏ��L�Һi):(EZ5��7T,�{��!�����OjƊ���!�A�,6&�sҿ���<$��ja鯆6��&֔U����B��7@=H���$`O�Ϙ����ָ=7d�t����q�^�IH>]�N���:�R<�M�;�����)��9�f���Ym�j�q����`-��H�K�c
��������tј+?Ii*�%��@45��9~���^D`�����px��0�q2e�p�t�7��=�E�lc	�<H�_����u<)&��.���~�Vt��}�����bV���<�́�(k��d�_���n���`[��(]m�=���A�=�n�$�%c�1����)�
ŞX"c��*�����*�*�ԏ ����z��ؗ��n0���?�C<���j_(Ӿ�e-Βw1U�1.�+�`��D�@��?>Կ�l��<Z�3>P����G�+�Iz)\L ��6�	^s\*t��b�4"�H�w�R���tQ1QxN�4�*v��z�	IC�\x��U.�u{ol��O��٭S��=ϋ+ut)���O^B��
|�I�E�afFY���7{��d}«��3~�����L����(�+}H�d���	}w��:E;�JR���[VBR��V�f�/�Ӫ�L� 7�1_CE�p��%KBܚ׏��9w
�D��.��銅��$G�w�oy�d����%��ϊr��2&��;a}X%�w�����.�zUD�4�����]ޣ+,��n�嵎"��Z��/���8��kP�yF�����z�z⪶��&.�#��3�	�0�Y���Q`p#��ϣ	F/��Gg�\��=�㶐{�A�ň���I�	��)C�6�ke��� ��*UU�v_{���
"C���K�)�@`�A��wUSJ�*�(<�)%�9����MWgc/?���쮙0�@�AF���͞�����h>��ۮ�ʃ�/D(n����:����W��WL@�ѕ���5�:�>��M�sV�g(�s�\�n�6E��;"��k-��s��]Q��?ٗٓ$#��^�_)wK�m�Gڂ��rpQ�?j-=���Q˵s��W�2�
Kԋ�B#RM�|�b�!�.e�kg^��`��	���NיB#yS.K �W�d ����z)f&���y�)T�����VB�_w�e0�Ć�\�4�3W���=[3x{ddOΓ^�I�P�H�ra�]L��h��,|ߤ�)�&i��v��Rg(�	��8h?����	�R�AdoA�� ��Wh�2}b��o3�d��1!pYj�>V����$׳�^3e�oƹ$�Uv��ZC��jDP4'���iCE.�S8X]s@��<7����D����\���
x��̕��T
J�_hh��D{��f ��ǥM����N�_��\�Am�U��>P؜���w��VU�E,�~��Mۍf���3�-�����L�*X�E�'Y	Z@���u�$�;��/��L]CF־�����[�u��m���AMbi6�/�pn"N�6v��E��2f�6�*�Փ�ک�!l��/'C}��j�	��%G�l1���+=sj���5��锝HϢ����J�f����4b.�� a�gӣֆE�S���d|�lSٛXcv��<H�!��|oD��I`��X�S�5�Q(H�tHKK�zǬ�w��s]NC��W|W)�U�ۑ{���\Kf,�	k�"�����t�*��
V�p�J���C�妒Z�#�Rtv�٠c%v�נ��м�_"�H���׃�z8V�H����Q}d��(N�\�{�E?{Z�2�8. ���y2�����YB��o��ZH�� <t.�~�$�U,��7�D�a���s����ƹat��an:���������И\/��7�}��uQ�&4	H?�t�p�]�C�[>+�oN�n/d	��K�;�m~ 46'.�&�֋�-��2�� ��?RT39E�Rh�<S'�V��o��侓�?�漏�Kܷz�A��r�~���h�$f�0"��Y]�}@f���C�TB�����Ʒ4f7��֞��DnYjz�}������1#�5AU3��D���w�hr�X�Ξ<�]��f�Iҧ�U�(Vy��۪�7q����>�D7�G��M�p���'��hYUw�]�>�O����L�4�=b�c�~O	�-B���m'�2��Hx֛�& L�*vo��\�A��n�|�
58m�Du���.�	A�߯��7#�j�P~��:C�%�:^�ZQ���Z����a�u�vnON��y��]��'���j߁4��ގA�����|���֫��׸b�UG�Λ�{���	�7�������Kn�Q���i߃┃���"R�[x�y^'�oG3�q~�(Z�K���d>��a�$�[9�C�/�7�;a?������{�rOu��o�sr���-b��K��������t̎K�� �������{�lS\�Dc�N=)�����)'���L�;�_Š� �b6�녭2Geؾ��`�d��nQZ��H�=�a)+���6�7�-��uv<G�u�
�}��h^0�+6`����z9���$*ߴ�M@
�7.����|�aX�_����I�����e8��~2���Mf�7�c%���`"�ʇ���>�ΫC�i�7�Y5V<�"�����g��������yYZE��� k��7rͳS�_7(S��m�U}���>��Pfz�!&4��4�8~(cA�y��n�������"�ۈ���c����U�����ٸ�F�l���YD�Dw+�TA��D���V�AXA7 ��Ƨmj}1�{�e&�����X���0�MB��У����4�j?O���Ў�p���������w��P���8 ,JKt[!���>��GO sGM[!`)�f��m��;*�=*.�`HZ8ќ��$J��q��t_!	y&���
� f@i�<8{�ھ��x����i��ߥ���k�g29��ǈZ�a�rZؘZ^��vϬ�J>�	ȿ�~D'z�D�
:��Z��-t��k���[Ғ��1��0�ڧt6q~x�2�D&�57�̝�zn���~D�P��_˽��3�'��"	g���z������&��l)e��Ht���IQ^׼� /�!S���.���� �� Or�����GC@��W�jP�N��)ELL�w���LxL�Ij;m�*Z�F��:�+OE��;�NI��2�x*��$4�i0J�5� QB�`�ֵxT�PuQE�Y:g�y�=:����g��,Y���SǱ�nԒtL!��˜,�2m���'N)�D�� ��sm�H�iYk^aY�[��5C����[t@��B*�Z�@�o��`Nŏ=�)|ᷴ���0Oy�<��,iN�吶(]��*�����龡�TpJ�(���o��4��̂C~��SX�Wb�*�s�!˛������~=��-O)aǰ*#�e1� #&�bvOVFZ��>rD&L����n,A��_xW�|�TŮ~���h�������XCV�֪.�'N
�	"�>����m���`Iא��)���6��0X�~?�e}VH�u����bV.�[�[p��s�Z��Y���aZ�@�<���R �R�I����[!r�o�6��[�!ʹ��h��k�L�&|]�o�򃥰�E:���p�~[z�t��U�%ߏ���?Z�k��fږ�%��T;�?�Eނ��������������������=������t�R�}�P8�����ۃb�{5�L���gZ6�0<���O7��S�M�M�٠����d��#m��3���;��Q=���=<����mk�hu^�����y�#u�;S�sZj��_}B���`j��/����P!VGդMe�>�)?�����/l�����ɏ?����gz�m_j�4�w��A�d]�;/� ��F{2}R��0D�H ��tV���gr!�(��XI"V�	O~o�l��S�-���-F��8�M%τ�#��e�]����}Ae4(x�B,<[%{�V��+�۹AH?�Q��]��t3�(��^_�v��݃��Eʕ�L�B��H_��	�����go֜ I<;��q.1�e1��ٜO5�
��|F�Z��i?wT!n�=no�Ta.dM
)���K�C�p`��e�R�rl,����k�S����<n��>ovW�-�p�q��ԍL�}� �"d-9dE�����x�UX����ev�J�ۘ�Ƥ��W���^-m�T��k��kAT���0�`7:B:���6����pB�!u����9� tbp� &�������Y&�Zd��*��㇖����nǄ!*8����s�*<_���g*���,��d�o�֥�k/�7Ͼ�
u]3�'��C0�� �٦k�-X���i� �q���b�w6[ϊ�,c*��O\<�3���')���j^��DB�>�ݍ�D�tj),�C/H2ؼ�7W�� �rq���g-�Xf{�4�-�Qu�m=�e(�
ܣ i������Ƕ��	��fၷ�������/���@���n��x�/4|�U �o��A?���׍�V�ʋ;�Θ=���Z�P�N���}��v崞E��XÐ=Ba�~.nt��`Q��-a�C~/���$B��`�|�a��&���g;�:/��,�4I5t8��`�~��9۴�-�C��|�"+&�&��z-5fOC�+��y�TX�>T�b�3ɓN`��\�H-SehS�5�q�־�"N��1�ɖ�B�D\�-���:������X;k��	Su\6�8qtI+ �촒�C��F~��m�R
	7y%�	E���H�14q�oJ�k"�S�2(W�${���m��l]A�c;ϒ��V���)PM���ڢ8���Y�GL�D�"-���|����F}6L�Z�i�$H7^B�9�������nk�)ȅ���ubp��Z�� l��3!�v�����#E���S�	����L؀�U������/<����m�c'1:�� �����5?�([O�^K(*��q�h!����W��c��O�ړ{L�v��M���Շ��0-K����T���40�2St���͎���9���U��j��۶V��?qѯG:*mN`qi d��ԋ��H���������n�|�"���G@�q�s����/uF��M�Z,�K�ܫ�� ]=�\Hy��O³/f�z���z v�W��t^�	ߩ#-jWH[F!�+��O��|5Go%�`����)��$3��ΈJV��q�Pҡi�4F���[��J��E*������YB��wG�W�O��7D����	41MMuo�F^&5�T��Z��HT6��������j�$�:�\#�J�QØ�?�1cyhXnI�\��{���M���($����2=;R����s�@�_������O����(�D�̷�b��I��乓8ܝ��.R����i�������J>��շ� �L���qs�N�?N���@�𽪘�/�mj,Wlw�O���1Ÿ�I݃r2:
ʈ�."Z�:�j�������/�0�'�m�Μ��(.����ڥOY|��k��P�Za����Z޼�!� � �ƊڅV��}:[�^��`�;�l#���$&�h��� �=$]���(k�fjV��H7�B���JX��C��=pXh�i���7��P�O~��|���lT��8�Sۭ_�Q�G1�F���3eB^)3��	WYa���I�1j:�� �$iA\���/�\ �JLl�\�v�{��S<���l�#���B�WQ�c�n�;��ۃ	�h�5�ڥ�,a+�Z:���-�,���;D�g8$����'�b�(�酯Vu�$ǰO�K�`	�f2�Ǎ��Y`�͏�z��NV����|� y�y�/4]��O'�~���[�m;[�eBt*��/��f�i��
�8���Q�����b<���`9y��&Y�p�7�Q����F|A?^�f<⃾�|�l?7�4߈��h�ō��Z��N�����n��0�=�D'Q+_�O<n҆��~O28_Si;��B��I�e [$�R�A��F5p��<o��D��X��P)���j�{���&l��&�/�A����x--�tCޘ�	̓��&@gQs�.��KGV����D��W�Wu����=�D_�HD�s�U"� +.���R=0�'�s�t#��d6���������cŲ?�H��&��ʁ���(�Ej����߫)�2?ujș�CF��z��������8N�._R>�@���nqQ��H<KG�(CLMg��������	^�����uXO�K 78P�9����>�9�0�D�G""�˰Q�Gy~��M^��=�E4��SVW(sqo&���iE��%p@���ߘ�7�&�hX�h���u�wKllN���M�b�c�Hm��6�3�۽�Nzz4H�#�\�ߖA�s2�t\����F�[\C�.\H;��Z"��F����}:D���p�J�k���A���nvL�6�t�]�Ҷs��y����/�)���`��v��r'kH
Y%��p*m݉c�p~�j�o\��Uִg.���6�sN����#F,S�*�4��[6�����ـi�
�}1u`(��`��.ͱY�99S$Ǉ�u,n?�Y�9�C&�{%�,���)�%i��&Q&/+:�93Y �ԓ�^Ã��G?3c6{/@'�If�}KT\��0؋���8�_�
��.��"�I\��>�V�n�u�%�17���_����-�[��j��W����d�Xx �	ۛE�Y���-ud0u;V�IX*퓌	�#���u�|h~~Ri�B��*àn`a~-�	lKR�QyU_H���ȹVT��Fk�]y��ʽ<me�����fߴ���Fe�x6Z�F�8e㿓t�Ѽ�5�<,Am6�5S�R�����n�$�l�����Ш
5�8�����V�s��-��S���Pԙ$Hdџ�VW����P���ڒ���U�J���� ���w��6����s�pǀ�>��4�ch��k�7��4N� +r�KI�� ��������'�N�8�� q�,Ϭ�u��m*��P�"�_��x�h|���%�¿~RiS�1�_��(���z�2�/����^J�?�(�n���	���V߻�Oܙ��'�C�@�M����2)ۦ�uٗ�<��9$�3�a��ζǡ�_̬�yX��-��KD,�Ox�QȒߺN���+�7�o���)|��S8���}qӨ�%�O�k��ٟ���&n��ot ˭�j������c%7��~�ۜ��{M�
��h�DF��d֕!ƤS��`l̫���7��M�e�ػ[��>��dlJ�zL�@��a�N#�T��Q�sB��]�Ku���h�0���u�
-����;;i�n0h]�B��+�˼,I|qb���ކ�0DX�f������S>d�u�-YC|J4I���*ת�������!�5�!~ނ������27��yh����Ћ���M^n�*d�@9�ӽ!:��c�ذW��=�_���ӭ�,�"m�j�ՔI�(�An�d��_I� d�<0��f�zz�5]7I�7�CSO�!��[��{�EZ��鑝��GN��y���:����O�G���hW\���@k��G7.��9�,y�9�f=��U�ù��@Cѝ�j���f�P����N��eR�H�$���r����y���4�Lՠ��O��5BR�a�.���=ӊ��}����Ԍ�sm����Kqc~��Xu^�D�L����!�� �_xG*�~&*��G��	�"xk9Iqss��eҌ�Z1_���u�����	���R�̄�]�>Ǽ���ˉR'��K ����=GF�k�м���u�ҕs�C5X�����F��hi���m�8�8���$0_�9���Cp[*�R���~�]�ݽ��Q���w�F�x����Cn�v�к�an��6�N�V&��]��4�,��
K(�]���g�
���YO�
X=�D��ج%H�����v��v!H\���:��^j~�Oz	?��-�΀.'��rZ铙PB��G
~-�0j���BȢ4s���܏8� *r'�M9����㪭�y� w^�(�E��o��bz[���i�c ��P��!;KV_�VA�$�u����6�C� �j'^� Ue�j�Hp�C�CrBiɑK��<~�XA���C/4e�T�U#�x�LK/���wPᄁ��:�H0rM���O^�_QA��v4A~Z���\�FG[�����Nv/0�[�-[�������,��k��f��X�[�Îr}��(����$�W����[�y�f�3����32�kfX�7f�3Ku���&&��W�I�V�������Z@.�7���m��^������x�p��(^-j3��C`@B���_��]3l9�E���6y�P�|����h{9x�?f�B%��L�Я/i+����j:N�}�}D��ץM���=���j��w�)8��#��u�/.��6���r��ո��-%����8�|�I"�N�XU�"Foj�r�:n�ޝ	d?�=��>�cD�C#;�@�{Eǘ}�*�s:��aZc�Z������6��V �Ej����Ɂ(����v���w��moY/ʜzm�bzyuΓ�B�/�Ұ�4���)6� WW�'˄ܙ �k���1a�s+��~�-?����C�� #T���jZO�۬�|ŭI��#�Gܯ�i� �r#�p�tc�i��_�B�|�ѷ���_Ӆ���������|�dHD#&5��;����o��c��7���]"gk
�KPH�q����*״$LⰍ��F��S��7��+��L3�@VBqE�%q�_s�i�A׵��$sDeJ�����B~� ��ku��T\�S�6R���O�q�h噓Ǎq`_p�Uű�l�Yv��1?�}P`^����!q�lk��0h�ȳ��T��C�rdL�U����X���e���v�+ȘMg�qs���b�#Q��F;�]�Kj俕.��`���KJ���� :�M�s��1u��ǂ�7-^;�J)��!���4�b׀���| �#=֚�=H3��4%�K3��q�b�����6���%��"�iS9�Td6�s��z#�e���h�of�W��`OS�o�e�W��$�!9O��]9�b�6f�f%F�� �#�f���Fo� }p�ss1m�q|Q�{�45�U��ba�/������(�\��Qo�����.;��Cxv'άH�.�����}A^ѐ@*0�Ć��HS1V�pΡ.��N��b7�gs?�2p�[x)[�a�@�r��}���2�|��eժ�/*��͔�l%����[̅�%^����ؠ��U�h��C4�P��=h��@�"3�@煙��jz�~��d�yr�=��2���ci��EW�q7=5Z�3AUQhO��o>]�s�;�W��'M\n��3Fd�W�ބ{���P����܆hT{���ֹ~���	L�z1l�nǞ����+I��K"R%�ʙOǽ7K"�Z�j���@*�%]G�9�9h���86��W��U�����y���C�<�Jn������{�N}]U5�k���n�@�.y5s��X��s�T�s�����v��SU�w� c,�4�6�f}j!f&)����]��ⶮG��d P?�ֳ�x�	�`����G��d�Y�A��������{I���SA�*1���k�� �\���<�|���'�2���ᓕ�^��ٳڬ#<~+3�[���y;�0�@��N������p�,7������{6��qF�jt6��L*�Ɵ��?��	�t��2h�h� �0�?��E�	ޒ(ǔ����X	��Gc�BKs{`�83�&.�ɣG���ng���c,]��3�;�&��pI/�l�B8�̕��:w0�����l��4�L����5u���ܖ$�M*�?�:\	���R{�@.iܠH��� �=�Q|���t�!��w�;��{_9���?�lW�V���}��c�L���7wd�������+�����?r��oJ��JK�:��P��j,�q�.�o��woc"d`Va�.��G����%5�8}��}D��_����Ĝt��&����
^����b�P?Sp��حU�H?�^���=a��?G�ya���T�[�)��+v������㜷e�yv����W�$��8�S����X	t�W@�8M'�C���Tsm@��%]�l#�h=jj���X�%�e3��BO�#d��K<�ig�g!N��7xN�T=�(e+'�x�llȵ�dWA&g��e����M=��ڛ�v(�|�@��ٿ�� ���f�9�lݱEH���]�vwժ��%�+Pԧ/ӟ�90�3^��,�s�N���J�dk�N� S�(?��@3?�� �y�^�~��`1��x�+�� ��>�@��
��Sp�H��Z�� �z�KNq��Z���"��i��/�򝎷CA`l_���ɶ�8����@�'|G>�x@�sf�@ü��R�E�s3y�a��u��*��} �2���E���]`��@��.[i�Z���i���t��[i@�3�,�ÐM��v��4��*�t����3��5X;��ˡ��q�64�)��	>/hy�ʩ}$��N��W��oOV���oCt�Kk�]/�Iꌻ���T��z��-��ĕ�*�e���CX�`���X���)O���fF����TjEZ��� /I"m�5��"�]�mpY�{����\��~q	�n�v�O�A>�!Țۛ��PD�7F��G�Жo)Sތ��~�~�>�W/d�,	0`�N|2Y�����4#,c��)6�yzI�r�����f@� U��Ƒc�{������|�gǽ$���ښJ��O%���A�W򀍥��e��`�u�`�_bx
mq�`����[e��e����g�gt�E}R��������4���[� �#�h4����wHj�G6��Q�%���!�e��u^���WőD�����յ�}x]���8Y��������yf�����%y:����c�ݗ��O�]�c~��>=r�xϤF�R�����[���a����?����l8��]{k����}Kz���|�����z�~��fS@���r+ݞ�lᗱ�ь�����$�<b��l����Ӕ��g7r��w'?35�0�/ᛐ��P�*yYs#�q	���Q��1���]mG�T���|LKЛku'眼D�[�BK
�_)�
й�_)Ơ$����8�	n�J��>�*�w�tX!� b��;����g�)��K�I�8��#}�C��dڻ�8������8F����zௌ�-\�E���譖1����T?'�R���0<�m�x�H֫_�;MI��E[ѐ�\+z����sQ�RC�%���ޛ��=c�]_�)�8�kw� |��P1���3W p���N1ޏ�k���-NLwx�m����]�o�x�w{�V�7�KDu^R���Z@��SW}����D�߄=r<��x�9y���,<�do���H��i����f�.h�]0q��4����9���NG�<6~ˁ�w�a���<��⌠��[��#��Ri�ڔ��dMI�j���p��Q
��7��cr56�uh�'mc;"�n1s�K�1���:�J�jM2�n���h٨xʜ����\h>�����6{}yu���i@�@m�#��,;�����NG�۳�����
�˓4c\�
����k�8<��V��5�c��4� F�R�h���7��k�X5���O5�|1I8ԇmٺ[����h|��.���L{٩�/�q ��x$k�)�ڷ�Gi_+�l�T;.�$��'x�Խ�	*[���̤����m�0F��2�.hx���s���X��6�uw@R��,�N>�A	�
.
��}u֗�fK[�}v��%B�W�e�|�e���
�v�m�	
{b������@T�C�Q+`��G۪Z�'����W'��b��e]�� �J������o�T��1�x�H%�E���`]��`M�34�l��h��cc[GB{�b��f�#sה@�+�݂/ S6hl��~��4��uUrM�8�_�C߱�R��ޮ���<:N��&Ѫ����D@��َB��HcT[��̳s�[a��%.�r9�U�*V�7��Il����pl��T��;� :s�-���I+�|��'���Q���� ����@�{ϸw�����d�˽X�Jl��&�W#x})�XG}���m�BF\�I?E����D�{A5��Q���D�Ř��5��N�
-�\��ç�e�7<#م@�و�SZ�_Ӏ���'-:��h杋"A5��hG3Z�����|ȑa���}_��ޯ�����"��^o��١��*m�x@�nĔ�'z�R��5�`�����&{���*��>���ok&��Lf��}Hԟ(Y���Gݫe�;N%`�9t)�޻���n!#��OH[�����69O��(>��0L�ȖA���)4|���l#FT\[@rD\��a��F���EPN��z�]�u�4a�{��9�o�^7�܌�SH|]O�a�l���08u9�Щ,��T�~7����६x�Gk�rE)���h����-9C�-ansn`d���p� :�\t�#�ܘ�b��PTA���m[r�CV0�Y���� MI���s�̑�r��`���6�T�X~��jК�o��������	������EY�M9��"�tϭ��4�Lc�J5����C��~�V�6�e���K6�t>G�2>��'��RG�B?,.�^��b���Y���;+G�_@8�4m|<U��ˮW��u�3�ٶ�a�@nb8��4�~�P~��/ē�ˬ�>�)���Y�މTӉ;2��2��[r4*�ȼ������C�'eprC,P��ީ�v�>���/pۂЋ�g�5)�Geii�Y-�
#�k;�`Q	��{��SU���r���eP:jRp)W�-Ē�!��a�%���.ع�e���Á��"|R�x�Q�q���.�U7>���^3Q$r+�ِ��y6r��#.��VI��J>��|����95�	!"cʸ��+��Nn#��WP��>��1qk��!���`�l��������*1�k�����Ǔ��=�]_��Ce.'D�K��t�j���&�@�e@"c���[h�z51�S�5��)�bqq��K�T���/�	=I�D82m�`�~M]���ZtQ�S�!�#�]�%���!��w�w{^i��t��F�\��J�ܚ��J{̋��.�eP�%6l���!���O�WcNb9�*a$��\�E�������;�|�1'ΥRp�.�>�X���~���W�����#��AS��F�f�z.����ד:����8Ż��8f$���[I�����0�xBZ ���@L�W�GO�-q�1�~0"8�{�:|�A34麫~�+\�]�f���D�|hվ�{�~C��P�=#t��N�f]D@���Zc��%[E"�����o�u�VI�V
8m�47�u'=.`���,�(�^��R��|蹗�}LV�����h���"�>�sy���K'��m.L�O�[u����T<j�rq���yIq��y�c��+��� O��^'l���+�-?ي:6]&��!�L�{�܉������}��� }�����9;�}'����q1o�l�`�XY��O�F&���f����J�<�</O�3(�o1Lc���(�����o�tN5����֍�+�o~����o���_l�<�(�����r�}dq������7�@J)6�%!	��5L��t"��E"QD��Ia��9#��D;F��y©:���7
i�ߢ�ny=��mD�oڭi�������9v��h�zB���/���q�A�Gp狡�9��EcMN�&���V��_%I����xD�:���ZU%ƒ����0˅6��nc�P�}k몦���C��Msw�U������>�t���,^�mH3��^�%P
�o��H�<�yet�6�,Eei&���t��U��!�4�[�m�8��ˀ�vmt�,��i�콶�ٜ&ܰ�S,a���ܰ�����=D�wS��;�]A	��R�,Kl:�:�j�!����!�h�����X��3�A��4��v�j��%�r�c�w���xx��{��U�C���b#��-Ӱ8���_�r8��7P�-�����CB�gf����5B�!�^�R]<9��碟G'�r�G��*�z�?��ѱ�.j�,t����nR�9>�yv"�&���^����Nv|-,u:|�A���Y����l�җ�4wɋ߽���Y�aD+܀�E\��)\|u��SR}P����l����Q.[i��F7�Yl�}ȲA/��M5ߙ s���b-q��g�#N/��'��N_��������r�U��e	~/@D$��/%��Я�)����@�l��=&l��^[0=�dBu����7�_5I�#P~/�� ì���RdF��]�jm2����I����8�ȺZa}t��1��\��.���C\���{���܆���z��p��DUA����%�#�R�3YC|r�By{s<{�J/�g>>E�B��
�:l�h��C��^��Zˇ����B�Fu��������[���&��z�	,����g�" tz�I��\�70�E����&!�� �6�V<�=~���<"x��E�Q�8C�q��.���������ѻ�MK���26 ���pMlW.tU�Lm�z��5�Fm��f�V�F�n�bl��KN�hbt!%�1�����ف⩭)�;�Y�7*LB]�Y���)�VV� �8$�,�!-8eˡ��m4��=�rR̬�4��C=y��*5��J���	͢!s˩�O{���h2�x����0CE�Ǧ�|���ӎ��}��>�s�bvUO�K��g:��H��G�.� �x�#�K�`���򠢧fx�:������,le���UUę�ܮ�=v@�&�CA��h		�ϼρ�x��fі"p���q��(��yR���2úͼp�c��O�y��#�ح#Ay�s��;A�}�4����\��\]�8��u��!�W�z���k���>
�0dx�j�gg�/�_��2���LO�'�@��PD�Js�f�&��f�������Դ�rg˹�sx��3�F���E�P"�0���J?�|�D��?T֑�M�C�W��|������ŀ��\��)�
����P�4z��+����Ɩm'��K�n��7�{o��!���p���"��r.���ע�D�҆��P�S����Y\#�������������JN����Q���4�<gb\��1��J�M��z�;��@��z��i�._�קo�[�'-���?�y�(EV�(ߺ�h��'�r�݂�F���sQ��u���(������?:�J)uc.�/}�>'�m7Y�c߽LK��_��pO2m��7��P��Q��P�ɍ%�v�cDV�WQ�B�v���?'V�RH�����Z��_Jhy}@�d/u)�p��M��cN3]ʝQ�G�u���nYt�ҡ?;,b��q��.pg>�w���W�E�I��2�of��]�H�Q(��Y�J<��t7���(��� ��V`��������*�ln�M4�30y�RD��>��^Ţ���6-��ӳ����[��p:t�^��(h�5
�����Ǖ=�"+=�M0ԯo�9'*��ԝ�s���ҳP�7��6bױ�n���"�D�Ȳ
%YsTH���[��tc�g��%f���8;��C]�P�s�;�țg���۪X���lF�XYn9F���ϓ1Ћ�5_.Qd��N�7���z/�c�6[F��ĉ�:�e� �4��h2�>�l���6$>� ���2S)m\}�&����^'FB��+oF�`.r<�YE��B2D���V�~t?fϴK�}�*��P3��C����pC&+�>�x�
��k}lAc1pc�z�Akt��%�-���u���7�έ]����ۏ���W�5	`�FoF�O��R{Η��\3$���68��ݜQl�vg����9*=�ؔY[�X���s���3���۬���0@�^˂�N*��h�5_���1'K�-kZ��j#ݒ�̬��D�x�3ܮ���;��L���w΅#��rν}h�vH�M
��)1sb\��k���0�Z��4.~�?^���E:SL���,��`����A�m�̜�J�*��>#x ��T	�y
�$��(��/w w�P4	,�Ë͜�VI�r���w����o5��(v�QM�9���η�]�)��6�?eO�*��?8rZvԆЕ�����h�(�qڹnU��c{�TYTQٺc�2��p9���5�%
ϙꌁ���o�i�A�������N&���qC0@���C�H/��U�U5�]��(�a:M%5I�S��{*���4H����`�3wiL/D߯�+K�؛�V���u%����2���Y�V8p+dZ���.�����t\/�����RX�1	���q;��}����9��PM�a�MӴ��7n�%��
 mY��T�5��P�6v?�*筤����lufj�4���n�ϓo��%�A��#	��\��mYG�#�v�N��N̛�@�~�CJ8��Ru���z�uq����*��n0��-���g-Q?Z��$�30�*��0�E��8���"R���E��8��d� 
q�tD�l�$���>14�xv	'~��Mo=͜U�� n�����yA�;
�Ĳ����b;o���	�:8(�涨�jP����"v�ڎN�\`DI����p4PC���4�yD�"�vjZ�6h{q:ٓP	��O�P#D'����]^R��w:�J�,��@�����qd���z�Y��wf�S:�s-
/r~{^YhO?u/��4Njlx��}�����u�Xۗ�|�\��=��%K�Czٳ���V��T�T�s9�<��: ��n;C!c�$�o�uMd��f�������;���o�D�"�5��Lύض�k��Z�&�F�'���sSL��5�[4O=o�3�G;��Y
�-��׷�(�e_N�B�MK9�}�a�XU�1�I���V<W-�QZ>VF��2m��Q�?����t�T����7%$lVJ�H��[׀ T�`̐����ZAZ����n"�m�4(^��Z܌Ez��4E��Y[�-	i��%]�'�o�
�X6��ǀ�3�k�&G�9�߯U����ŋ�ڍ��I҅�^��2K�+����`�?Ix	�X]�wk���,5��n?�e(LQ�v��7�8��]O�'H��.ߒ8Ť2���ݘ�]�F0���8�CEN Py�6���"96	%��Z����uC��Υj�;��X��3W6e��Ƃt�4���nPTt�F�U*���t�	?���5+�Du�I�won�\���z���I_��ҷ�������ɹj��[�>iOC��z@1�J��U�TR��Yg����pP�{��@ξ$�5J� ���Mρ�œ��)ؙ3>���F/�3TU�v���8�FV��������Z�T�u�����-~�A���()pDBd�)���12N��A6���)y��]������m�V�t	lB\t{�\��Q~�.�3�"���\4�	El�e�d��^�DZ�&��,��{\�J����&F��G?ͨ
�|T|mlj� ����=" sͷ��lJ�|��8#���N��oذ�����N[��p��z�V����!�VE
�×������sv��7($l��3Rt7\ϙ�H9%*>�Cu����Ul�8 ��;��^=�Ś�s���� �R��qfAꫨ�9b1@�!3��mk�Y��������歅V=�������NJq��u��V޴d�+3�s,�^���}J�C2�@�4����̵�Oٿ��E��0uV�[�F�쨿J�����������G�+�Z� Q�T��r����������w>G��w��V���mb���S��TM�w��8�9���V�e�g��y�rm���Jo�c(���������2����͎�K�A��Xk�3 )f������HdPu�(vL��:|5�q宎��|ۜ!��Hc6��N6t&ŌX�c]�w\�<:�yT�e����h,BH#=��d2a7S<�g��X����(���I����
��ĉ8H�?�q�x�#)��]�Nz������ǁ���s.��[��K	m��Ϊe�Z������#
GJ8g�H�M��_[ �������/��:�9�wf=�aa�G�R�H��иj?��p/�
%�'�zu�-��殕긣�nl<��������&��s�V���S�6�)�x)
R�W�r����� O^�S�g3E����ΐ�٣��c2����˶l��,�-vr\�r$+5����(����J���ǩ�@)�Kp�I4�� )�ӿ����w?ق���y����
�ٴ(O��s��|�-Jd�jO��L��P�@�x�7̱r�{�D#ѝbs��e�	L��nN:����ϑ���@z��O:(Y���z�	��|�J�!�zJyh+y>4��'-t�����v����Ӽ7B��2RF78��(������*�����|�q(���]�Ċn^��`'����vI�<
�D�x�f�R5`8n����W�$�V���f���J�|,zD�N��d���R���Y5a(`�SgP{!'��.?���]�o^W�9"�����a֟��F�(m�k?�^�%V�8�3`7���Y����bhȲ)������[`
�;�1u�f�6�����Y�L(q߼uz}�h��9����Qyhގb�a��<ER�J2BqG�VRK�(�iZ�z�R��%��h��W?���������[<ˈ$$�[w��<+��_��vXR3���IB�3�Û�B��=C{'A%�<�����9O�x�S���[ր
^)]D���y�+΂�L��m��D`?B5ׂ��(�N*X�TX�
���6>��j&{��ї�h^�Zc	2t��m�ř�,������X'AZ�?|R��(J�^�ˈ�+M� ��%�\Ұ�@���el^��7�N��%TZ�mv���_(���̂�u(�r����HqK�/\�
' ��3δ��y[Key��s�a^���sM
�j�\�����:�]7�ȍ�$��'��Ō����0㌺*q��ZE��@n?�Θ�fT�]�rq���nI��b)(y�X�&���r�lA��9�������w%��Ղ^~��W)嚑
�|P�2��	�X��)���ۻ}�7�Us�}!��y��#HC�^�������wώ���Z����=<��5 ��@��J[�Lx�I~�@��%>�����Z��U	q���
8�C��Pc[�l9֖s���47�˻0TY+�}�{F-��C�4I����t���lB? ��R��菅z���7;2%��x�gx�6>m����Ah���A`�&�L񇆰My��ɡ�v����@� ^i4���S>Ċ�?��.G��H�z_�e��#YBh�\`Eu��C��t*��hkAo�B ���z ��*�Vn6��S��c[���<�C�H��#~�r?+�
>ٲ]�ϫ�:�:iǍʓ��df��2�w�W�? hm�������Oe�^I;�kH�d�@R���[��0C������ɭY���O����/����g���+�٣&Q�B�`�N5��N�����ɼ�R4�4��
�eg��>׶jO6�1�R�:��s���K�jyp2���9'���S��=A�A�u�Lϣ ��5��p(Z��&������Cd���������)��b�l�.��϶))>X��K���	�ܾ5���
jS����2Y2-4S��u�1~ '2�ߞc�RR���2��o��B����$��������k�d8��/�RQ{� %��N�����E֭���	�XR�k�|��K��%T%�Stz:Qf���:����K"��`[*�k���WH �91��Ug��*�b'�?���u+����5��X���εt(��N�o���ezK�H����iP��@�P�29��O��{3�i)H;����W���x�'�M�<�Y���\0n�P���y�1H����Ӡ�R�Ū4R�ߝѸ�]Nc�^x�;"4c��K�tڿ���|�O�P9e�M�yԨ����Ϛ
0 ^)(��bJ���[���*�}'_��Z���`3�$�״+���-Y�K�h�=8�L]W���T���W=ݖH���V(���]��C��
����Tt��0��>M�ۄ��ZN�] ,fhA������%�59�B?-W< ��Xx��^�v�.
��E����چ.ڇKB�7w��`��zS]��6��'�/�f�)���7e�}p�g
G��5u�����t�mCb�	��?��e�K�g�Þ� >/ ����C'��[�6�q����9���L�x+z���>���l�{�o�Ї��oF���2Rm�cv��ۺ���(a"�r=q/z�<x#l��J��Sgm�>I|��ϟ�,;�]��w_<x�x���Z�?���m�	y���߻�S����U�O+��f>��g��i�l z�1�$_n���:"���뮲�1)�"M��~�s8UW�bu����: s�JcH���(��CA
��=RΎ��,1Q�iy��A����T���fDɫ`���\I-Ϣ=*�?MLPF�Tei$j��f�u���c�o[�I��]o$I4�姃^ ���h��p�[�����K�e� eN�;��S�v��Б�ئBL9'�	b�b�Pk�3�G������6[1��C9�v.*������^�����"!�ڽ�+�G,������ioZs������F~���Q�3�51�Si�!>�V��J� �%�hf"K�i慳��z�O�f���u�;Tg����V�܁cK�aRjb~���6��Ƙ���9�^v��2:�� 5�u���&
@U�c}x@�>DJU�Y�n�X��VzP-_;;V��w���s]�|���ɬ�^`@��/���@B��wE���Blf ��k�Z!(�C"*�$�Lç7�B�.�$�M�l�����I���iU�q.��&��`�������"n�q�\\c��0�etyc_�f�;ᮐ$ópC�q����!]���e���ڌ�+(� 	�=-�6F�<�z��>Tbڥ���>�2�Zk�P�����w=~���o���a��� T��Wg,�A
�S�	x`~�{,0}�>}4W����Z���QV�C⯁�|�c���c�c��9�.KЏ�/��ï��z2i��/���`��3k�:/`�=�zA�#������En3�ߠg�/�j]*I,�	E��t=�u�3Y��}����s�+��c���� ڭzlI���0Rcv�$�X��[�+ƌ��C�	6��%�"{���q<�����b��Y�j�2����Z��~z�X8� ͧ�%L8>A���!�	�IB�[K2����x�Fm��E-[z ���M�FжLn0?�:�N�E�^F�
�������H)�����R�+p|�7*��֏W
��fȒ۫�_z<a
:n;�*�(C��3m��.#�
�AFO�`^��.�I�����@?�6���Q�MR��d��|;�+J���5JE��?l�&,D��ҭK��W�f\}tf?͝՞p��4����i�s��*��V\.:����V2Yje��臎����ԏ��"G�%j��Fz#S>�%p�3�
���u��7��B��
���z�Xb,u��=�c�[���AO�eG��5aeto6���C��S@h��z��{,�L_�#�<b��(==Y��|�(}�h�h�%�!����k\�?8e��[���N�&~��&�C�4��xOQ�H���!��g��r��g�[�P�1A�,w_^��Q�}OD�<i_�F���z���7�3N�������.�<���	>�P�L2�� y��������s'O���K�o6�͉E{�	�,�F{� ��ѫ	�BL�~z�݇~y�w���J<a�6U��P�N����P�|�+H�`
a�Z��׿�һ�bHY������	o�78FU��n�u�z�9�v�nժ�ֲ4X�_�2�Kː���?>�|��I{z�N��Q5�o���x�P�9����q��>��t�Ge-pO�k��B_��Y�jL-^{@��j�qh��Rn@`Eű�v��Q�r2��`fc�C�c��Z�%��6�z�'��T�dOS�7�F�W�J�;�3���"��:b�G��
V �[�H��A�)rR�#L �݋1g�E��M^R���Ie��Y��Q!xW)q�����H����0m��)t�;Ih��|�Y��/d�õ�`-��_Fz�?�Uw���mM�mJ��4�|��ԦZ+K}����ma}�jܶ��,V�L�5v�@�#�دG�t���Xc�@����aL1c�WT��n��~/J+pۄ�-�l�J:��󄧗�o����(�C����EzX'D�-�K���3Qd��;A���*�t(�c+����ɓ��Q{�$�d�ov�'�W�����p~�}��Vb�L��EA��,��d�$��$�;O�Iީs@�:�V��M�х�,L��q�7辩�B����%������r�������G�k	e��?Ѥ���	("o3�� �I������L]�:��EY��Oƴ�!Mр�!��d�9e[8�,|�r(0P�h?뻈1H�u��1(����p��/�`���d��:�O���k�buqg����A��Ғ�d���N�]o������)F�xdX��*�*s^��^׻JɄ��{@c�yK�FNۃ����U@��y��-��≷�jP"m���j�Q�K	�fV8�B� C����d�Y��B� 3�(��#�i1�����Ҷn��B��)��>o�*�F�#��̇��1{��q��Kb�P{��A���axk�Y$.��Sf$ӳ�%��`�>;B�����Fy����0���Jл��WO��*H����+���:)2�iӓ&�Ѫ2���?nq�Ƨ�sX�ս��Bьz���/�뽂��9�B�l�� ���"��61r6�g��Å�E�Դ)@�a�'c��<V�_w��˯I-�F7h��iZ�<#��`IpΔ*WK���PQ�0�/8ʥ�@4�@����1|}0�`ry���g}P��VV)3��R;;_h�_p���Kjwɺ�c�~�v��w��i����~�j���u�$k�/��)��7p��v~��:%Dil�p�]��C�*�g�"y��[���s�DqK{	/7�Z�C���(^������d!��5v�nr�W��\�]
6s�v����
]\�m�P�?/:8����v7����.�.�M�4��`�g������m����6���y?�Y3I�TR13���O�buW�.%P��UG�WhR��i��n'�ʍjrS�J��I��
1�5�����utٍ7I��M��WG4�	BU�C~n4ul�&���LW����"���h�Y����o"Ӣ�K���d��;���o�#�Po�7ɠ��������{^6T��F��i��d����}d��Q��3�ˢKn��j��l�;���L?+NC�	2;Mh��@�\�s=��]�Yϝ�v޼���؎�p��� ���	�d-k���i	c���p��U�� ��q����@C��,`Ұ��ˢ��xaSX͎dl�%�V V*�D�;��8���}y:��A�؝N�Hj�p��}�-D`s�W��;���+�Ӫ�Q��)�2*���؂zY4���@��3�Y�ϟyr.V����l��|�~��XM�+��T����A���Oz�lb(ZP����c�Lhӊ��5o#w���M���K��v.M�/"�k�!Eu�nѩ��w���(N�B�Լ˫���~y�k�"����D' 3��k�Y�L��fs?2�NM���sS[�~��a�g�u4��*F1�P?b��Y�X��	�Ӎop����B�	N���Q��+�Kd̈́Z�U�/HC�E���:����5��Wv��I��G'-��+Tf'�tY?�3:N���S�������?r7��F�0�����ĺ��mK�2�Z#|���"�D)t��D��o�$D�8ƤDΣ���O;Hi�c��g��X�}w`�,�}��
��HxPϞV}��g��I����U@%�_�.Iv��*��3A{1�n��81�;��^�YD�p��.A��c�[��O��#+%�Dҭ����\��!��]W"�����hse*��,ea�4ͣq�7e����}��N�y6�jK�x��!�� z��E��(���V�Ӧ F�\���׍���E
#�/S�Rh�9�s�O�5a]�e����led��{I���}��+B�~/�B�a�=,�Vx����������hz��v�@�L\��з��jX��Q�0`�x+�r1��/�yE�F
n�@�l�T$�c-` �?V%L@�D#5:T��}**i��PoV!,9k�c6�+|����kݯg�#Z.{�nƲw$:Y�P �=t,��?�M)�~��QI����Ɣ�R���RN�jS������03���Q�Yq�̽t3L0���w���1�{h�Q+�&6Z���
�6�g5��[tz?��J]D���7�P�#|���BY�@�ֺ |+�m�@0�@��gwD�U?=�-���Pz}P1�iQ��$�0ʰ��D��M���"�Ёd��W�7ϱq�2�;�Ud���˺�`�4"q�9��7�h�_�۹��bZ-͈ɖ꽻2�T>p�$'}��E)縐�$� 5��O??�R1��R����	4�t%ݽ><���*I6�n��}g :0�K��p�]�Ij� ����Ҹ�^e�� ��V%�,���s��F��X�rt��_]��G��.kG����^�҇� .Hu./�P.�P�:{��ܗ�g��ȁr���A9��.��g��z�c uG�XǞ ��|�w_Ï���e��v�=d�W]����N���������?l���9�ӵCU�Ɇ�L5�
|Wo�1�}e���+Jn���N����y��S�
h(:}:<�`!�y�fNG���Və�JGf'd�X�d1yqiHuH��'C���IS�̖`s�0^���^t��:�+���W��ڒ�X[?�%��r���/����T���q�le&+c@�Y�q4�^��Q@*}�6a��"@mMj�O�[�t�����ݞ�-K���x
k��:y��x��,�|_�7m7�v���� v�q,5K�2�L�s������DI�1`;Cgޭ�29������K+	�{�[C �E2ࡹ�41~������,�=��s<ڭ.pH陣������o�H�ߩ��"o���Sz�3|�8W��t�A�x8wҿ�����3œX��ݰ�ިйE���f�W��lx��p}�p�F����+$���Y�?$��/�w��>����������t�|k0��T����5�<�l�=Ԭr:�W�#,����=��{��yf�soc��'���3�	_~h�x��.�`)�.{F�~�军�q'�f��֏�O�F5�bƺV�qN��5D�� �&A@
nAt>����u�7��D����T��5z�<&�>�~G��X��:�"�	�>-"Ϲ�͟k��Js]#'�B��y�sE �wo7e��
i��u++52�e0h�����_<t.�8�^��.>]V7���y�k03�.�{�~%فE�)f�w����F�9D��w����ç�6�y~�RȀ_d,�����R�-g ����&�Y����oAֱ�>�UB��S'-�����`�nr�S�A?�O%�5�>4��/��1$�H:@+��Z�ĪT$&0bFgW��cq��ɚ�5�%��r��O����qC�o}1�N~��d�Q|�d��
���\� ��Q.q"�<�;��2p�S9�p[ T�v��Z��CwJQ�,ӯ�؉�U��$mn#4g�(�{C�`�'L\�gć�U�> �C,�[��/00K�_����Z��aR<��l��zi�1���
�`��E����3��-�ޛ���
<�ko�p��}ϯ($�Z�X8�nC�c��]͜~�	~T�6S�T[;RY؏����ƪ��g@~,G�@A3P���R��]��`E$v����0���{�?�%�༷�K�����|�w��m:J6�62��0�j0��z{�r�����r����:=+��Е�Yv��m�훓y�-'h����b-�����R8G�����"��Ֆ	�J6��)��z��%���p���r��,[p�UG2�:���~`M��R�m�4�AT�FT�M){�)�5�*�J^U��=��K��e!�1EM1�6�_ #����)�=A�h:��к��G��E�&O��b�Զ7!�G���f��0j#I��>�P3�k��d����w�jE+䳃/����i�"ּ��&��{��?���/���|�e������mck_�S> �Lb뙺��69��by���ѱ�D�)�A���+RW���ڶܺި��B�3hC����2�T�P�L��i���\,���u��$�HxEpF�7~�s�A�kWin	�(����;Q�^��������v�Ү�su���lE�:����.�I!H���ڻ�ئ^@
C��R��G�_U��|640O��gT�ʵA�|г���������=)��k*�j�<H�c�3"L�v����?�Q�=�K@$�[�׼�J*�m���%>�e ׆����#ޢ����c�f���^�m1oX\�4�G>~T5@V���{��̵�y+�G�3�H���������+�]��$��K���0�)F"�n��s�/���n-��NH�})��2�<�ᥕ�V��}8��A�)��/5S�߷�[0v���07��[�F�f ���יB����+ �w�\��%���$h�c�Kl,���$�cc:�݄���x5��rY{q �T5�:�#�%��x�F <�%���gQD���J ��b�e��\5U�M����f�높�O@zB0��m�����������-ʂ��[���3��X2?�Lb�
��?�m[����E/~1�U�
9�
�/HDf9p=�ʩ���@/��".P�Ț�������"�nl�[
J�B�T_u��B�E�Կ�FS
Y:7���mWO�ڿ�{S���l�ݯoPR��x>�%��jwGb��-^1�3���k���t۹%�01�-�IΩ��)VB��S9#�}�b�!���1�+_�����������kH����z�CQ�X��!�,��37Ӟ�"*� C�@��Խl�_Щ@��'e=���t��wx=�`T����͔��@;,K6d�-����+[��|��f��V�����<��xN����G�$�U5KA�Y�3���m1z<j�Xc��1�?1��]ʛfޞ,?A������
p�*%�X����.kM�Ա��*/����� �4_�>�4\~��P���_�i�a�����#;�Ab�k�����2j��<�m�t)_{������}�c�����t���1�ټ��4�:����B�l�|s��d��ć��JF�#�_s� E�*�(YH>Gj�Ah '*}L���И�Q�\�f�.��$l��56�?I�i�7ixY�3أ;��UIx˒����OB�)T8�,�\I�
|���J@��W5���̵��pw.۞�� �p+lR�D*��"M�������m8L�����B���P'���nʐ�����*#��JB�	��0�x�_�}��p�ԅ_�μ�S�7�!}��(;�%/�����$8S�&�m�;�r|���sS��5��K��/���O��<G4�Pv=J늓V#��`�4Gq��A�:@X���rk��pB�,�~�J���uC=q��;nЅ���J�{�4I$��pYI��Pd�/�1N�U����N0��Z�������8�d��l4�1�)��gX*$(� �5J���F����x�) Fb�&LU� ��/n��lnҫ�x�a� #C� ����LH"X�/���'��Zĉ��Kێ�?�_ʹ_L5������C�1ɴ��C㮲퀠u���+�f�v!���Xu�hIkRٛ���K����;pq۠�B�+*.���.�S�I�c�PM������ �6m��!�I����׈2(�[={�y+i�\��Q?��a\p��-Ih�(����ßc�^�7�X��9L��C���@^o�Sh,�1I�~T�M�Wuv����%�A`��{(��E��J�Y�N�85$#�eG��B� ɔ����Wm�QVX�h�W�"a�rre���)�K;LA��VӜ��yb����`k��~�۬��ꞤHN����|V���k1�eݽ��N���e^�\���zg����֥��(�x2 ĖHYM�Ր���o�2��=�fh��0d�$k�ewC��9<MP=���ia��/�X��9FF�����ɋ(�8�7��}'?��� �Z:m��� �EŊ����\qիUԄM�Ț�)5�ӗ�_��4�g�����X�{�W�ygĬ�S���r�K"�u�7	��b#9)�6Y2�[��vL�ނI+]��ߋK����V��3��{�(�~���^��	mrc����l����un���қ�5Z |��7���p�	T��'�=Y3!S���<	~���j�$*v��-�c�F����G+�r��[p,��pW���D��N[51�>������1�d�қzs�������S�����ùԮ�o���Vd��k6��7h��3@<�'U��t&�|��V�H��y��M"��+6��`,|�)RH��_��_W2@��j���m�4�i��IsJ������o���(�p[G���N�< �i��b%�d�T�¦T�<��9�4�]V�`b�w�W����Д�ν/:�}V�j<˙pS#��x@$���H;��s��l�.���/���`v&��t
K;�f�_��{�X�\)����	�5q?T�',K����!Nxv+�ɡ���t��uf��]s��Ie�����:2� e��Jk|��]��#	�����m��M�oth~�����'���?�)XvſJd'�b2p�R�WS�m�~�pj�P��}u�������e����՞���� y����D��չZ�@'���e������_M@�F��|��'���"ё�u�Ac6�Q����4�A�
��ZC���F��� a���D)���R�^m�o!����*�o���P�Sv�3������D����3�C���G��OE �#k+Y�^k����Σ�l>���
��t��:c�����a?�R-��P��&D�K>*o�Ǹru��rL6}Ƭ�N���d:�0���	�fέ��|�/���fë��<׾L��#�u���u'��_�j��9X0�� P&F���;�H���W��:�}B�[d� p�o�"�Di�:ŭFpS���~1�21m:��K�绷�U��2��Ra�l�7�o.�bDy�l�@S���HNș�#��S��6���;5{�'-ER�WU���B��s"�C��,g�8{[��5LO\U�9Ɠ*�&�qL�x+f��Q�+CA�l�R�;\�:��~$�Q�6Z�Yc���Ȭ��ܸJsM��Y9k,���5ڨ�ufIr'�!}SP����vdVk�yֻ�UQ�����Iu{Yc�R^G�-�o�9t�Ϊ���㱪>�ľ����������A}++�܆ 5Τ���GY������A�#o��G��fc
uL�=�kT�p��Zy�֋E˸��TM9��@��Za�z���Z�B.ύ$���;AOu;O
�d"�l��.�����������ƤA�.�2��N~ܓ��*�ێJ�km��t�1�'�h�p��;Y�cvZ��)发ݸUt�H���b��:`Y�bdn�z��a^F4qX�[g�-�^|���sL�T��9�+��U;���Ǚ�����N���vZ�Հ��K��7�����>0Mb�1(��~������}�$�mW�-{�@�^mˊsD#�Ǭ"#��wsT"mQ�]!��l5D^�=1�^��=����Bn<����� �ܮ%V^ȳ�]�/�}����`�#XgU��ƪKl�����.h3��aH��wlZ("�(�%	q�C��/�Q�(?�٥�j�H���ކF�������ǜк�
R�BB��X�g��y^� �}��%��MY<����Q17��0 4s�~1���~e8.�ؖ5�_:s��ʛ�YE�'�"�FYan�틯V�  ��RK�`�Rŉ�F����zR�1�Lc���uN��ߦ�c��=~�
P��cD�2y��L�R2�)i�G#m�3�+�l'�{�W�oo-� R�(P���g]2�qu/���٨H�
y4&�����EL
�7&P஀�w��t5ɷ�$wɟ�����%��S�46�*-�cV���Ή
���<1���.��V�tIK#��Q\����j�G��6(ƛ�9�����L�L�O�Z�ɤ����s��8��A�b�����@��_^�z�t�|�Ȫǩ?��{VR����6y�"�L�H0*B�B(:Q��˫��~>�7�z�yh�9�����J��ށ�e �����F��߅������Fу=p�0��cW�'֞�����g�^�j��Yq{�=��U��V�Z࢚l7M�돁��{�[[V;#NF�����J��� $��]R�� �(�I���'�8�sϧ}�Ny!�xF�Z`�K�� ��/�l�򉽼�~$��*�{H&U�����z��i�b����O`"Sƻ�At2��'d��㥅�nJ����[��e�MT[\�p�m�u��P�
���0<��lWf[�a����=)��p��xo���j�g>l��)�h��=N|(���FgZ"�l�(B T˕�G�m��PU�2D�j��Ǹ4J����#n�.�V+��Z�ᆾ�ͣ,�w�u~�S���̥�ؙ�G�d�x��0�r�,�P�Xw�S4���$�=�ΐ�C)��!*K 38�7��Q�bE1&�Y�{��F�"�^�]��Y�=�IO��~@�
$3C��'Q���}h�e��`\�L�IM� ����`;���o�����%&�����a���}��,�1E�V!�7M+~�ج�s��� �zQ$6��IV�ܓ��rj2����~�hb�'��D��^� �k0ٴ��v�Ā�0�D�5�T7"������б��~�ci����X��Am��&.��j�Y"�ʒ����B~��3_��=�M[�;�C8�F!�hj�x��U�ȧ�m�D�W��#�Aw���(����}FpUL-Έ���c�����ꨱu�6�q�6��2f�-N�SF�,��sM_��γj�����X�w��Jcq�"˾ً�4?��Ͷ놛~��v�C�Ò���o�z6C�p-����~�c�F'gaR���U>!�&�2A�Kq�G��O�avH{y��n�(�Q�D�sQǮ���{9mךL��vf"񶅓�!I,��d�gf#��h����W&��C�%+��z��\�wQķy�Oq��v�2$�����m�k�UV�b&� 0���{�T6Γ�L�4B��I/�\����c.�q�6|H߀n�8����4�.C�	+.�М�ULY3�(ik�=R���s����� ��t�>�e�}$�6꫟�!���A\N��7B73�)V������E��724*�����ӽ)�cHI3̯�?�JcC;�!�	Ѱ�0�#_~����<B�s� jHG��'Z,j��k�r�hڇe��ؿ��n���f6|� �r'��s	��-�c'i�FβM��v�,�m�k���1v��v�L��;j�
�y�����xQSj��!��T;hqa	] ��m@�7g�gg��@�`t�����YoGT��ƛ�/6��;��u���n��HQjNd�A�qh]��Qu��f�P�,k�^~)��KW�@�NiPא���"��׬��Ü�á͗o��D>Dx$U���9d�T�s/֐��"s���;����E�V%�����+��07��J��YL$�+-\�&k9~�VG��9�b�zX�D��]m�v�?F$�ыX�UŇ�!-}��+�P�W[�|����$�n�6�p��_�p����{���e-c�َ�S�3L��<���u�7R���3��H��*�g}Q���2�bc��k�/��R�dT�a�a�Ad�J����u�������7gtZ.eF�fHT���G�l<�{E�Զ�\�֟�w�bg;s��l��M�Bq/�r�S�m��2)"p�Y�A?���>j��O(���j"L�잮Xgx7�=
�C0��S2�\'
�e5xy�R��`V�؟�MwcU[�K�K1�B�a����k�k��	1@a�Cl�M
'�*�Qy��ׂ��m P桪�%��LE�b=Uy1X��B�ڪY.��?<���f����TlQo�R �$�����2G�[_9��+�Zγ��zi֟�.ݦ��
B��k�L�#���5q׸��F��<�6	`����=� ��}�'��GO �s>(z�/+�\D�qJ��f��1��p��)��?t�	�ҕ}���r���H�q���1�T����G��Qz4#�����L"�d)�[�w$N�L<�O���%�}s#��LQ�2�8E=���<�+�N���@�9�<��27tI��/})���P]ǎ��]2�+s�	��7�7>�!���z��wP�w\�v����v*h����Kx�	��:�o�����#Y�SҰ���Ү#���/���7Cf��g�P36�Qk�w�t�b��1D�xsA��I�g䄝���>D�,|��ĕ�z�,�	�$���� �Z����cY*�9�72�p� �5,��{�\gN2A�g���<�Þ���Q��-ܴ��tglM�n�uh�i#O�v/��U��C�Ņ��B!r"�򊯿�.Q-l���� �vkY;ƿ���j�(�ڢ)K��3{Ñ��VD��[�K1VJ�����+�m�4nS�+�3[�������Z
F�ԛ�g�ski�Z<�:�&�)�oMМJ��c��Fۏ��xi~��.)Ӊ��>�b	�1����z,m����[[>�gH�נ ١���-�G4ڲ�2��8�w�w����ɵ#�TO-�<����a�����{�:pd������;'����0���y��h7z�g����q�-���8튍<D����}��4.�*<*p��G��ΠZ	^�_񉀕J�:�O�)��XnU i=� 7#m�v~���[%�]�D��op��s�/��}����9�ƄM3���u�D�`u�&l"ܕx�`��S���=�\��R������라cv�K�q�;|`-/��m����|���"ƥ?��vBv�����p��r���a�2�J���A��\���}f����C�=��o՛v�һ#�{Sتf�i��k�oOpIW�H����{�VZ,���+��ڈ[E�{��o��9S�YѦ����BT��m�=+/ryw�� �g����}�0W~�3 �+��cg��p��q��7�E��N,|��z�;a�1�C|�1mX| ��&���e�q�uټT�_�G������m�0�E:Z#ٻ;IƠ��W<�u�G�B��Z :Ok"�g�O�n��Y�ƹ���D��(鷔z��\h�t��B�3�HiwBRשyX�H�J�s��ʿ<?5��u
bؒ���
Ȗ0�o<�n��w��I���LY5����߿j�Y�9=�SPI�C��;�>S�����������O�r�cFqƏj�e�%��3�`�:3��ǲ{�J7�1��5�7w΅x|�=���?�=/�I�+S�^�X��_�6�+P�KnyڋcDf���{$�2(ݽ�\����g�-7�['F~J{H�n�C�ۤ�t�𷴗�))��%z���~��ۈ���,�Uܯ���ĕ���7X ��fm�u���f���{���N�Bbb��ߵW��$��o���4E8qK���I�I�ʤ`Q�� zlX�?M!�Ala@`�����Ю���w4������e�$��|D�	9�P����:�Y}�Q/Y���i�����M�-��r(=�=Ҫ�kM��%5C��h��V[�ԑ����ŉ�]%Rw��Hpi�oA~dv������U�UbnE(��`�s��^��VEn� �t��*�ݥ-*!`P{�rdLH�����$m�Yd.(T樑}�Za�����5��w�V��W��i���S���4�q^*�Pc��H. ۠�~c��$~/�U^���KK�,��3�b>���O�p�^~�Q��*E�1��q�}�¸['9|��WTb��tY��#����ݏY���U��]���	K������)@`�S�\U�C�Z�� ��oa��>ͥ/yP@��
G+f�h^�G�o��J��甘5�jkI0�I=���J�5P�ʄ����ג�b����}n��'���:T;b�$ȅ"t��GKG����*�ӒD��Y���?�?J��*$���&�r�ۯ��p�A@1]����z����9,����ۏr��k�����'}�z�Ň�����d�ȋ|{{뚟̒4� ډ�ꝸ�q�1�m~Z=	�n�jAgtEB��.�7I�%xr�8�_%�Y�=�_�Y%r[��Z��8��������3���{s��u0;}�T�����-���I,!�ꃏ�y]�l�uۄ�3NO�2]���A��Lw�o,��$j&p��YW&HM6L���[9����WԒ���_�zj�1?V-��ge�SRYB��ṗ����E گk�27�QϜ��uH�P��6�d)��o��4��^���=Z�k=��a�d���;ԣ)Tq��I0�����"{�\t[j#�\[K�V`]!!N���y�U$�^��xF]8�J�lƃ倫>�*H���X�;�E���"��+��.;�p�+���g�!�陾I���������C��ۦ�j�/G���1���c�൞ڞtZJ���,>�[(0�^	#K��"��
����;��=F{U�#��LO�c]��Գ�T�P�8_"?��V�Zsކ�d�IN��	�+�^�O���!�D`5�;��ڑ�8)�ʡ����M]T�w?N4�,٫/£܀��6�,��'���J}���e��[�Q�W8���J$��U��Y�n����)��B�6���4X8D�f�qtc�gS�mv�l��˘��H�	wV?�� ��>84�cC8␿i8�r��ܠ�5���+UX"X9��S�<*y}�G6�]s���Ag@	� �n���1����5��s矇J!��G^����FQ;���>#��W�����f�u���c���?-��Ӻ��b�KO�
S�Z0<hř[&���^r�X���dT��r��S��{b/)��qF����!��4{º�?M�L[���^�U��^�u!uȧ�vvO�� F�����EA/��$�2�<���Q�8��:����\66���>{LN���*�b�A�~x�<�`�P\@�eO��Y�y̺�i�qi�*ΣV���o�t���[w㓊Cχ��+�2�3ʵ�w���P2/���Q�x�?t�c��-c�ւ������Fal����+��Qk�9-�]� �}(I��qS��T*h,�KO�8*�j��f��E^ x���%�*�bƂ���f����#���_�5hڲ�T��,Z����D��O��k�{/FP)��=%@Ή�#>b|Ri�#Έ��g#c��w^�ou;۸�%۵1K4��73��o]ׅnG+R�@� k������sT\A^�Kؕ�`;qxpQh�����3Z��8
ؘ�k?kL���Y��B5��k�nS+������ �uhU���ģ�g��|`�Y����O�����Y䣘���궘a?��d�"���y�V�:� ��*�Bړg�d�'�g��q�U�٧���<BS��(�q+�ﳴn�op�G�������y(UѰ��x��yb���x��FrY��[+�4��x�C`��a�!ѣ������^}�q�^���O �ݍ���v�'V1H1��L�r�=|�m$���9�Q<e)Y��K�Y�S*�u���%�s�ҷ�-��I���� ������j�$�_���*�Ч�e��BU���~4�P�����κ��nY�=3CH@����Q�]�d�����s�t���E�&�n����}�D�4j��'����-˾ֶJ�'�v��TN��ZiCBcŚ� ]�{�/���25��\�s�?M�&�~;�����v�P&�P� ����z,��8��u������`g(5Y�1)q�\~�|� э������%!s4L���O'>7���غtOC�}���o���f�~I����#.8�����:��o\4�zTɑ��H9(t��G�A�lǒ�.Q���4Yr�_P��|D��5�)�'5`��N�I�Hm��r3ֈK���L�~©<S��8��߾����ȼ�X��^��<Qo?Z��Q8P]G��d#�0�Mk�X8����d�`P{�+�+,���8�n"�Wۈfk\��`<�Zj�J�HїQ���Y���y���4%L���q��Y�T՗4i2d�%PB^J�5/<c�&�y�*�n��<����&��Fdd�{p&��b���Ҳx<�zbf�ٍ���m�@@����;�Ԫ+��,�>���6O�җE�;�� G�O87�ә��B0�K�% �+�P�Ę2w�S�K/���o���.��^�f\^}=&�"�=��US�����˝��%`�;�|�*B�:I,����������h`1Q��V٠�/��(�����!��]'2&�O[�:/�m�%�l���j����̠�\+�8NA�s-g+�d��e�Iװ���k0]�e�_+�_��1+�E�J�b #p3�.����r[�����p;$�(p���|{U�G�YP^�Rqkj(��,�H�C���Ͽ���qnD�(�6!�	���^,e�bz]E�(x��k��� R�7ִa�j��=�Wd��u�X'×�h�ۭ2��wQc�4�|�.茪��8?w����PO�Ĝ&w���Q�%~y\�]e�~�a�`���q�iN�L[�Vz��N��I��x�-�3J"~�nV��c��N��lU 	?������Z7�|E�b.؍�<x�
�k�CR�ѵ�|\�\E����x]���1-�g�K �:���=X7�q��)~��<�úw{Ή2� ��X����ϫ�]�j)z�L7��Q�Ņ�`ˤ!��O��,7]�b�ϥ� jy�����R��<�;_@����E�7�:��ܜ���i-��1<	l�BbM�3���p��z��vւ�[�*�Wߐ4�E�D$�
S���C%��ck[~�����8��R�;��)�휵hXC��|�yU�0S!����Le�z
Z1 �du�����>]���h8O�Z\��E���j`���o��^gEF�;��$����R��@���F���ǎ���4Y��S�]FGډ4�����>�$ek�#�����6����c�]'�}=z9p���21�����QB��⡗T&3>�����L�����������S�`@bQNg�p9��f%��d�w��_
�ML*��[����g'�|��+~���f:A���ՠh�E���T��N�;�,'ǘT ��7�s�#���)Ȭ
Q�+c���S�&v�V�n*��@"b�u�P]	 �R���T�K�=��~�����A޵��y�"?�!V���6�	 K�P4�!�T�V��T�2��a~v��V�E>�ߏ�LJ�ž�� �0���'�f��nZ�4⅏�ƹ�=]r`��K��!�V'��ˬ����׬@���U������$^�P��?#���сn�]�F�%R���1T�l^�+/Mڄ94��i[������|d��A�������3�ǘ�4z�%���O߸l�O�T���Ht����&��i����t1�@,dD	-�○"��M�p���G�b��kc�Nx�b���,,��5.�/vմVE���ڣ >U��{��u͋D��RD<����]���o��P�7-|~�O%���ɚ"tU�H�?G`��I���O�_�Q����"�%���� �[璬�L-9P~���!�>&��&v��嘀[�{�1�����cP������4�zDW �x���V�7�+j�\b��(����M�3�XĚ��4[�8Yk��\πW�I8�}6E$sKh�>FY���D�o �ߚ������p�k9�=�{�1	�gY����Bۛk��P#M2��F��\'�N�`p��0
��s�}/-c�
w�J���D4��z6=��%��O�j_���_��w�q�U�~sf.�4&U�C�R��=ѷ$����$ړ�G6H�"����+U�ub R���u�1Rב��	#��B[.v�5�*�4�뱤}M[@r <ͳ'�j':�v����c��~'1�Ym�;�)�x	�dX�`�F���O;cb}���9L"d�ʗ�#\�"�skjJ&����������jm�e�hS���41g�!�	�5+���ll�	����b�Y7u٢��O�ن�}U�j8-�C��P$�b\��^��&��$��e��l��P��\uD�����(;s2��'����r�XE�ƥ#WF�Z�E�`I^�8l�R���j�ߍ��G�V8`b��v	�+�ȴg�U ��AJc�G�Zό�WU�{і�C_hœ_�ج�G�}G��J��u�ˆ@�����*G�ݘ�~��S`���s�����t��SE��b���u� Q��x�GF�����t���&�L�H&s딭��]M�����C�z��+b���Z*����w����׋�w��!"��F��*
�W�����+%��M����D�l2�����P5ޏ���p�Wh%̓���1�BhA��dQ]�`�"p��n}�:�,�]��o�U4�Ba*���L<Բ�#8U�3�a=��+;�ƙ,��=�Ӱ�����^PG�Y[t�,�`a3
��_Gڸ����x����v��Q�G��<Ԉ��Е\����S팈i/2z2�\���ц_��`}1,��#���D�JB�G�%��P�A�6�_l��Go�F�M����<��� `��T|<�ߥj�ۛz��'O�H%>|�d�@)غr�)��@���B������^�X���_���[P�|�|��~=u��/�<y��w�|�+*s��ڪ�&�?fn�l/��Bġ�R[�r���4&,@�)���Aon2�p�#�?�.4ӏ}�����R�^�|�(s�s7���9�<���Z��Uzߖ�
:�'KO�+h �+|�������NH��Q6���Z��n��~�o�g��^�� ����#e�Q*�������FB\=9Uio��4�I����q�}�&�B7غ_�8���IC�5����$�4��F�=z"��'�z�?��t6~�1T��h�_E�!h�xV��l��rV���'8�-Y�i"��Y��(��Q?#�-��Q�TÙ�qjyTH���L����l<h}c������
]lcq�O&�1ܓ���&6���]��`%w3]U���&CJ�i왏�����(O A���aFv�ܔ�'M��B�Q�eR�Rl��/�h���%環�� �y�SG��Q�u xL}2��ҫ��k�k�X\�JI�W��y���E��q`���׃���MC�;*^�p�@���ń������t��(��/h��u�hG�o^.�Qc<�� 3���[6ӟ�<6ߘMS	C�WĲ��?�Te���l�t�F4�� ��;��6��u7~��NG�����z�!��~��W��L������|�E�+{��F�� ��ᣉP��<2k��pzr��FQ�`�0���-6��&�dgBQ����5(.J�t$ԝښXy��n�Z-�����h��(��� &�a���Ƞ��TU�;Co�N�	� ��k���E	��X��v�"��~'6I����d.�rgՀ�f1�ꂞ=�����N�|EUܿ��~+����vh�~JͤR�D_7
oг�N��̞��|�۩���s$8bS�D��È�>�j�[]�1F��ˌ�r��7Osi���r���I8ۺN�¤�.��v>/�[*��4�[��h8���J�q��3��,��
���%�;<qI�#kU������q����t:�¯<�a�:te�G��k�k��.��(�m�xs}uFJR�d�D���#��Zx6��t�P����F��b����K�m�x�[�89I���(S��'�!��ѫ	%���m�)��|��-�%[�9M�O^x������V�}>t�羋C���ő�����?���#��qp��	ny����gf�7��+��< F�y���*�ۙ�N��d����Jyo_,�n�
����v��i0�+��m����}ͷ��qp�\��ZƧ���S�q���!R�E�7;^�SA�iHs:᝔� ^���Y��c���V���O�(���t �IH�;�D����?ҭ*@S��5�O��� ���'Z~��I�1E�y+*�r	��bF*�oE��y��&�?��A�<+�1P��S��*n:�Q�[����P^��:X
[�1W��Krǃ��=�d���.C�ZL�s�W�!��M$����]��(����S	�ZTt�)߾��r �*Fl�¼�rYvq=f�k���)���&��ni�d���k�e:e�(/�?m���qZL.��KO�����ϰ�����]Ɂ͋/%�ߪ ���Şb��#1�"�?�j+�5-]�/����:��|�!<"�3�U����'�f�ڄ?'f��L������0D�~třJ�JF���.P#N(�����x��Z,/�pm�ư.w�ElGD�Lv�ZT"�9�i��LX�����	S.������H����?(e:1bqd
�$��˜$&ʧ�*K�-<۳�Ix���a\$��܎Ab�u*Ԧ��vt��̂���h�L�}�%�Q�$��Ӳk�Ϸ�c��)�/qޅ���@��N��^�F6��F����Qg��-URL��|�nKr�5[/f�/_��8y"z��@�5s+����N���Vn�Ώ;m�T �=`)��1�}y�f�I�\Eۮ' oȟW��z+��֝nl0GFe`��?mn����S��2ԭS����Z�2_fذ��!k��Y���G,���ߧ.4��V��|M�4�`�=���H��Lj$�߁���b��)?/�݊q����G��9�,5HnR7ޏ�~�H�vE���3Z���2�_�(+�i��0`w.��O�
1\BD�[�7`��Q}l/�tcg;�����D^�d:l�D��ˣ�й�@�p�zs/̮�Z�y5���B�fs�H�7kB\������F�f����'?/�HkA�-�~Ru�-��@��t�jWc�ΙE��x��"��N��C�z��v��]����ӣjp	:4K�[ʏ%��KG�G¤�����k*�Ht.J78��λy\-��Ėq)��(�E���fS<x��I�r��đ$�t~����8�����5���,q��:-m�� j�՚y�s�s9���G�s�p���P�R*��N�k�Z4�^nA��}���,��^��^3i����ǟoz �#��[�y�k�9~��T}�w���3���-� ��=�k��C���7�N �ІKp��)�K'rqX�DN��c?�� 0b6 $\.2KAQV��H��G�HP�_��F�1��p9��fK+�MћIu78�I���J'��{V� ׋ًq�J�������߅n_�Ǻ�;@Į
ǪqZ�ѽ�g�aJ-UB��Ѫ@q��o�)O_��O6P1����q�Cxޚ��3�b[�B�:���|֙����j���}'}ΞJ�!๏�A�x@A��\}��y� -`�V�h�y��~�Ƹ�ړ�?���P��GZ�TK�|ps2䟉ZL�f��\�
�B�H 7��'�a�D�e�,F�Í��ub@���J��T,˃��&ӜdY7<�\K��(�!GW�x���Cg���Jx�SӸ����-Ɛ%9�w��lV���E�����;L��pI�����s��g��V�������M�j�PTt��H8K��J�����z����a����F6���?ϝ���l��^�2�/��1Q�H��)���]g��!�t��͓���h(+|[��І�07������]���63�%(A�h������eu����%'+1d�����	U�7_��1�ɪ�v��E?u(Ou�md��|�b��^�~��!L��F�>�
_ҔG������c�$M fɹ��a��j2{r_�.@����"s��ͩ��ހ����?��O��EF��Y�y1����Q"r֙�b2(�Q����.�>�&�na1`�n�f������W�77�v��Wz�b�1��8ݡ:�~CL&,�!DI`�u������Vu�Lue�[�*�w��Ga�Z&5�?�{Ն��+6���{z�_��������u�8<T�a�羍�Z4V�m=J��-�����K�܍#�7��ғe��L�_��t�yC���oאy�n�b���<�,��!:ɋ2tCl�L�3�ĭm}�����J����q��%�<�Oz٦ɎA`խ�_kJw���9hw��}�AR%W(4W�H��>�G�J#]E5�{1�u�.��]����Mu�\�[1c
�Wj�֋�u������E
���M�;� ��is��-�x�+�8��T�lё��N'�{��P��am	:
M#��z�KC��ʈ豑�oC�>�F ෫�׺_h!n*w���猑��'[	��ٛՎ2D�?LJ�4 ��Q(�tH�nȸ� )��|$W_ �n�4���<����6����+~{B�V���%˟ZMw������k?RV��4��Sŗ��������=^1�<��qm׈ߌU `�;����\U+a��<�W���W�����h��&�hY)���S��Сz�����XR�g�+U�l�y�EO��YdW:y��]��t�b.��r�.f	��.�⭳ɧ��=ԇ�eeX��^m�(.��!��]��=�U%��N�d�%�J����4vt`j�R�J�tg�q�#�hHC�RTX��v��
^�]�Q����1,Ԁ8,��>����u.<��K�����ع����UF�~/�Dq�ЁE���IDqQdp"�{*�\���\$[g��մ�q �%�2���Rr���P���5������	�U#��$	qo��`�B�ƘkLD9L����=1�mERxJ�D��s �?��9�\��/�V�3�FE��b"%���`G��oХ\�� ���h�lX��ٺ��F�����N��):���7�=�1��T �g?����8����,cs�����t%߷�G����LxX�;<�pT�G5�b"ϱ�ny/��5"���>q�߸���F�R�-�g��l<E|�po ��w�)5{�n�+�I��0����y��X$r|�f%;5ڢ�JQr�-���(6�9��k����e ftb��>��ZqBY�JM�b]g�W��>2���+W�߳>����{�����_6�_q���K&{y�;i������՚&���%�5$KR���$w�0ck�J��D��
xa0X7xWU�����gك��W�3�s2� $�`�����J��%I���ލ>��d�*��Q�-F�$V��0X0�;Z��r� �=�����\����o޴�,�`)T`p��f���rNvҚm��iZ�[@ ��H��%f��в��܃�䪝�6\ޭ��ߞ#2*{+MƾV�����
���j
(P�H*j7��t֌K��r$��!���J�)��.0BN��pK��_x��|C�U�H]Ƥd R55�����%?Z�~��f�S���N��y�2N�P�%��r��"b��}?{*o��p=�_�jQ�JY���.4� ޵2}̻݋+��g�7�KM���F4�����,5y�X�8��K�a�4|�h[85wE��jG�zpie��
#�~�G:�d�Y|����'���M�ԉ�E+��9�����v���>T�غc$�>*�@��Kj;�Jr��4<����i��� M_�*a�f�|���-E��s׍[��ds�{p���7OI�^=A!M�E�?]58�������^�,��	��UU��B���=�nC���BŹB��eD�����M|���cac="�͢�\�so�~D?��	�(�@p�IQӯ�8�/����WJɉ�Bf?�  W�Zg'n3eէT����Xs\�����w�2BczF?�T�˱��f�>�BkX�{N���Jg�2�M�[t��FF	5�a�k����q>�\���JƜ���:��M�]�F�-MQ�><c�*d��mw�uR��cu��[�}+�ٷ��b�vј�Z���F�G�_m��K���fA�X�w��/Ϯvg�O*��&z%����%��s�6e3j{TtҒ�6�'�����ũ��N4�0����;[ղ�쟆�飺/��mv/\3��K�h cX _�Hp�J���}AC
*�{)O�ئ�2PN�]�[��X��%�Ϣ��0E6!n."��,���5����Km�y�m��\��_�� (&(:��f!1���>���a<�H��7kN�۶p��;��)��"16��v��# S���@f3©6���b�"�s��\rS����DN�ɸ��[=�fpןy-���gE�������['{F�;S7�|]�z��x(vFB{0�Ԙ�ԏ��Dޣ��g��u�5�����%��y[x3{G~���tӛ�D�';����h���2�F���ר�v9�WR���!m��t&	L���G@;n�ٌ�1&ұO��\�0��QG� ��<a�x�����X�[ӮkHMj��i 6�d�FvZ$��V2�k�]#��?,�|9d!��\��>���P]��|���gS��$���Ŏ9u�(�8�n�X�(��񟠲��h/��K�� �]F霚(��\���L�}4[!���o�es�4����>�#Ay��	8Q6����%��ȟ�ZC2`"8�.`^,�jgn�,::�&���*�s ~���������뺵��@*'b��Fv�;�x@=�VW�6�LL�g� Nã[�æ�V���w�GEw��T"ב��"!�ӝ��!�칼�x؍3B͞r�OZX���J�V�
�WQ�f����oF����F���������rkO�b5Ż�'��#��?�f��R��j��`yЖ%\�t�ۧ���q-�N	5�շ�W��4��q��w����%�du~Q�ozG>���]�^������~�3������;�pjiO���	k=��?���!#ݗ�%�'�KO�z$�0���Ͽ���A�i�i 3 �뭬����,<��X���;��!��R��n�Ti�f[D-KruCP�)��@��m>hH��U���8�GxN3�f�k��u$(�>蠏�����x�^b�!��I��g���f�ң|���-j�/C�T{���}S��۩��Hi�`+,�T��p�o�v�������GǄ�P|Ȝf�4D0�ٿ>3�-����׋�À�V��!t��ީ"m`�3��ȄV`���0�!-�mK�����|e� ��˓=S��:M~Ly��(��N�=7��e�"+�\��}J�����
�Yb ���l�ƜoU�08v�>#�����h_�qL�SUL�o
>��4���'�d�2���݌���E�&�[�v��O���@j�/f�ն�}ӛݤ$�Z�:-X!l����Llfݳ�	���<�V7�6$Z.��P?���	R�ml�>4�107Z�i}A���gZ_^;���@"?s�^\Ӣ��]��0�j^B?C��kt��N���:-e@��a�r|_X�ə̕����6�>]��瘠�8��z�W���<9�hQ��Ze��#_�|~%��Իu�p�He��y����"0yNwǔ��-��O�ƴ,Τ��r^�AşÊ���yŠ<1eɓ���TG��^��Ɏ�_�����J0��9��06e�Q��B��{�.�{�������|@�b��h���Fʐ���w���$�YYU�~�ͺ$w@�RHd�s�nR��4�p^5�(���?�+䒶�>�X�j�S�3S���8�x�\���*� ��T�:s�N�� %�)�J�MF4�طȜdW��t���v:JAK���]����N'ǖ�`��=����.;�ô�Wz@@|��3��&�pH)����������4��X�6�����������>�|���V���#�� ��H�>J�����wmyV�S����x��I��O#�����Q��}%>��U��U\�#=T$�dF��E�@�e����a��&ƽv��ç��p
���j���į,o\S�1���s׈�U����	: ��[\�eˇ�� ~s��I�/{��B��n�}A��G20(����Pn�.�~����Mo���}�V�g$�&��k��� �]@�Ǧ������a0�c�`���(���4��a��8��ѿw�����7Л�(��$��g�1~���9�> �q8
���Uhƿ̸��	�XN0�0M��/
�{�#*�s���Q1dj@6n�Ia�CZ��n̆m���id �Gd��c�U�(L��⴨9��W]47|�F��)f��fd�=��&���D5ڣ�C��{����Wdpk0�	����k� 밋c�)�꽑�.�c$hEM��YE���z������t8<���ŃA;���1چժ��pF�9�����)��ظ,,��� ��{����j�0�zuX{��a�W~ �C���|�FVZ�]d��OG�h���Z�6W|�hn(��8�qT+!(�'ϒ ;;��8|�6���m�b�-��/ʟ�k ��EaE�W�N���BKL���ReޟR����f�"4���N?i����p���U�A�A����N(���α���+sԾ4h�9_�Ac�����ڞ*d��<��\�v+ W�|/�Yt���WHob���҃p�r��\nQ��ծ��� h��E�/�J���2�$��������%�J	M��g�ߓ W�)��qy��:.���l�S��|��ҵ���r�Wu1�~�/��nmʅ���0ޔ��Q��U�k_��Z�:�"�C�{��)!t�+u4:���L�m�3���lp!����d�'�I�;_��+hm1P�;�(�j#�2�:��C-T�[sy�����c|��k��t�l�������Թ7�aFG����p��`T����HԓU��[��#�]��֢Wr���%����[����-wV�V�}b'fH:� ������E,"�_|�oF;;!"j����5���骳���p�<�ؼ���9��Q ���#&�Va!�e��[����(c����gb����g��������@>(��pŞ�K9����x�p3�p�����~C��,k�u�CT����'��5�&�w"
�����4�oN��	����
G^ǃ�[<�48?�CW�yE�K���`z�	��`�<tE�oKa��'��{�I���И+��}��I}���2���<4�4�9m��O�0p�Dj�?AZ�s�[�3۬�*JN���ᙢ���k�՗�0�W\w�h��)H��V��V�>}�9�Fð
�c����|C�%�;hn]4��Ȭqg�K�m��������p<���E!����߅�J%۾�#�5#G�~�H��D�)?W�p��1�PT7"�)���V�	 ��É^�L��W��;n,�,`���o[p��uuc�+K�DU�e���e��rk����vlS���o�`IU��VU�M�m�r�o�+h���n�9ƽ��ѝ���j*11gs�`Vw�(Q��V��Y��C,��i��	��-"�\H�9�S��/n�Xt[���%<���~�O��x��x��bZI�~X���3�>l�<`f��s�
)i� U7�����t���ԗ�JljD��x;�Z �_ެ+�F\�n֘����$��iaQ���r$�V���2Е�-��H���r!ZޯI���j"��M��ػ���#�<}��/ɒ�T���C�~V�(
a�MܬCOn�������@�tgI���%��k�{����mSd.4����^2�3�~&��>^Q$%�^�K�h�Y-O�'/���_��z���;�`�ຨ�D����Q蜘QVX�&�5����S�kMG^�\H`��	���&�{��W���F��n	3�C����C�ަ�eG;x̷Odo#*5!��ɿ�h:j=�a���}���,�	��ÞIQ��h�yD��:u�{�MУ�:�/h1R�:��ܧ)pܻ��I���u��R{����r L�ֹA+��b2�LO�Z7�U�:�|��ulM�k��QI�4(ϠI���H`�3�w��wk���J��<O1T(���_Yu�?�__��d��.ܚ?l���M͋8w;��}!�\8]��-�N"�,r�3���}�v��j�rm�a�)�0�`����*��T���֬�������M\�8�6 ��*-@�} Լr*��'�5Y(��6��L��n�sFҀUP���Ĝ$��ڭ����2��7�~���F���9g+���Z�����\�n�E��Y�����cb6�y�~nb|���@�a����E��s`�)D�\9��i	�7���*�I~�L|4W�D�*��k��ӯZ$_=�~q8��]l;�f4tH]�u����:3.����*)ﶽ���M� '�,��9�`ض��8+J(U���h��#mӻ�c8{:ȥ��9R�����%�V���=N�*�m;l�F��L:vX��l�T�M��� 8�o�Z҂%7��Vڵٗ���Yjf��Ԝ3����å��U���9N_*N~)�*E�Y�+k�oˣe�A����ۍUrb/��.}~�����'�7��v
�:(�
�RNj�"M�'����y�.($��@�)�<��y�d��W��
h�I���9�
���PiR{�������L��`q����U]bn+g�b�QL9���6�d|�Ao��1鶡봧ȼ�Ì.z��������+��m/�����3���`����ǔ���f�K�����L�t��H1�)j�k�L�=tx2b�T�aX�F��ZO�g3W�CVq:�*aS�G=������	Z��I�D��o����Â-v��:'��x�9Σ@�9Y,MP���1���=yu�{%J��	�-`�{����~ׯ��N�]%��^���V-��n$���ð#��T�c3���pٱ��@9���D/*F�>�ӛ���'
��D�?�	���43m�F����>��1�[c��,>ӣp���H�I4�BM��>�|? ��L��݅��8S�$�F��SC��G"�f=�g���z���s�LE�0�� �@�1��i�H�v�HG4��J������\�3a��]��:Ľ<�p3t����^�v�Fy����g�#(#I���T��'�T��.����S��$���Q���̍2���g�>��V�K����V�PԁY˂& ��SD�;֬ 2����S^'J��Bb�T���dj�bK�	Y��p�Wm�Xg���T$�bc��3L{m���_v�H"�����ӺN�R	�c��	gh��";3�`���Z&�b6%&��I��ֳ}��5��ڔ��0������f�Oh#����ԺQ}��JgN�@*=�ƴH^._)>�̹���Q�C7^��.i�#�c�@M �K����������f��K��H5��%�?7B\�ީ_���
Uc����N�\Z����VL`�i9X`��gJL�XߦX��b�B��u��<���:|�DR}yE�({+�umΛ(�SZl���q���D��)��Kx����/�\l"r5�fK�g�B�7@�
*��:(<���T��hn��\PM�.�vj��?�O/���� N��.��U�ߵ_Ȓ�����p���cup���Ђx<���^� _������X`�I�#XVlD�Ơ�����	�ĭ`�;�����s���IݓY�J����4���3\��i�ud���r܋��/4s�﭅.���i���<����O`M1��L�?�ީ]��w�}w�h҈m�#Ԡ@�YWcߌ�F�4n�6uh��M�t�B�_�B��{E��N�����o�2�Z5y�������c���$������#Q�+j=|�^sR�ʻ>�M�M�5�[=,p������w2S�۟���ED̀e��mA������1H/�c�O�=p�W��6o��@�!����	]=�����n�w���?M�gJD^oTd8����k�ez��V�Q<Y*;���+�[US�����	֚B�/ۚ]�\L�%��	��co3�Ĝ��K��Dk:ג"����ߥ��΀�>$x\3�R@��� 6�玞�mK��d%��O�F��C*�	o�f����#"�
[��i��ȉ� ������ܽ�����^��P<�?�P橝�~�xS�����=~C���*�\� x-�ʆ���+YJ�g/�� ,�n+h�g[�_T�`��\��\
P	jY�|��6�IҺ0��R��Q���C����q������!	�S[,����H=b(�c�sl�NS�?�N�L����0��C���*:�xZ��M���e�-��^����_�ʙ�;1</�۽"Z��-�>ͥ�s�h��K���r�>@�t��H�u�n��+��T�Dza�>����W�p�:iL��7�^:�S�"bE	�q�U��x�-�},�Fs/�+_��wޞ���Q�y��"`a�dpA�*,B�gM��E�7�E!(ťD6�����G���m�+\v� �R����"�h1t��BjL���7��}��Et�T�ҭ��_9N6'n�p^��G�lXk2����G�`tV�7z��}��n�m��
6ރv⽭p�C��b`e�1ߐr�kcʣ�׼y7��h]t��9����lv�Yz��!�!E�|��f�q��[�m�m���P	�ͦ������ԮYC8�0�(ݬ**"���j�B��uziO{�;0���~���FQN�3�O5�9�$󻘴�-�o$�
�i�R�|KdzS��fRK�\9�t��O�l����~�2���w���s�!?{WJ�ӡ|Ҩ�.��$l yO܇]S��ю=H�|-�_.�䲝�&�� H~����uoF�Eu�K�rd��2��Ќ^��T)e�DtC~����b�!B�g��]ƹ���6id\"{s3�o�yA�֗���=�-���)�Z�	G�=�G�٪�`A�L-���MVw�2i�-�q���5��J)q \G��-$�:,ZK\�Ғ�B�l�in���s��۩�|���ʲm�E'��`�Ի�i�`$�Ȥ�WF��]@aШ���H���w��J���u?$wD�I�I�=��G���ϡ�m�aj
��3�ĸ�ɴ��a�[�996H��5�+	��?�=V�ez.���&ٮ|����>�K�84����a�0��Ů�T��Ur�}¯���o367���1ʔ��1��X��x�c3~^�cFǥ�ξ��a�%�4'<�^ߊ��� s������۬�������#��y�zdA�]��5���_��ʵ��Q��ڣX��v�����U��,n���a�n�hRK酙�A�p^�g�ZWqx�c��<}Z��� �V�tB4�1�0��s�:fS�LT�_h�X�r����6cnz�X����[u��-�l��f[���#��+�"��;{l�"�@��'�\��r���z/m,�iE�K�|��@�)�f�gs\/:1]:L�P��#�&��Qf��g�w�����F]�����~��f�#�jj[x���+�����$�u�Z��T�¦���=^��2����:үj��+D3nB�|�j_7�6}��(ٽKp5��&�.v��N����l�J|�X�<Q�JD��-�� Q���O�Q��$I$�KUV�͕ #�B�����8��'g�IZϹ�������j����!�'h�{|f��]�+�h(^`N����Zr�YPK�-�	����*��Y�H/���^��>�P��T5$����ʻ<_�r�L��(�����&DI$}PH�$ d�/$d�(��S����t�ѱ\Z���;�	4(R�^�S�0yC޹b%�ݘ
W�`�(m�RN�K(v˜��	k&�.P߁40}�L&&y���RJ��9�J���ʝ�J~U�f���h�̩"�O��gȗ�="��s��$�����Օ�.�n5����΍�+W����<nS��֢���ܯ�zz-�3W��-K�Ag�bD72|�_F]�O�����K�E�;�Ƚ��[�de��1h$w�I�7 �O_��h�p�#T�)�	z���CC��:#��800���<b\�~~%=�����k��sE]q��-LT�u�p�&S1�%a@��=�l�+,N���j_
����io��nQ�uY<��v�I��Z���\��%��w4痰Չ��n��Š���ػ'J����0�W��"�B�Ôe��s�u2b�V�Y7R>�o, ��z�a��h��K'\��V$'�]���qև��R��z>	���~+͂�����ݼ�>�m��?Jj/���Ӈt	�E-�m�ۄ�������`7�s�=B�9��p�ǿ��� wJ-N��4@׃��9���@/po��/`8)W�H�%�W�*�����W,mv�Xea[������M�RW"WnP���2������k�#Q�����=q.���ZK�)�ULvb���t!o3M��_�H�R\h�������Pa�k�֚QQ������08�촛��գ̓�0���+�,C���!CG�9�)AW|���Kd������G���O��F�X�hP��P��/�St+��Y�E���x���_O��*%z��T'�m��¹k �&]�:����F��>~{W�����/��B���z,�w`��C�&X��� ��#�֤
_���olx���Oz�..�����HL[�ej�=��C�2y�cݼ�>nȖ[Dd���+�ӥ)��ԁLH���]�ldJ�?��3�'k��� �F`� ���áЫm.������%��(��
Ti�;g��cG�.����O��zC2�=P�~��L�@Dc���q��"�@�G�n���:�jb�ѧ,�J�tӋɮ��;������M��G͛��hӓ�kPՠ���ȿ/<�ƢߍV���o�WCA����'|�e:��G��n��_R��ņ����)n��0>��ۡ���*t�|��й	JH��?
�)%m�*��#|��4R��C`�X�h���)G��cz>���{}���j&���乄��PQ�t�6���Y�6��R���:�� ��5�����"�]��ph!�Y�f��x!�+b��0(	)��]�U�0�6%ae�܁����4�?GF@E��Ƶb{r�F�$��Y���SąӚ�Hҡ��P���Y,�ll�5꾌>r�1so���m졦����1�L��V�ŀPx�e��H�����I����΃���(i��H�F��҂=��%��Ò�vf�E׮�Fyh�T���*e��;�(���q��H �k�F�8���[}��n���(m=�Yl��S��Uqb�n�OZ�74vH:��1P�i��i84!Ya'wY�O�uH��z�Fᐪ~#׽�I�5�|R��{�H�����d��a_F��َ��ko�٠Y����Uq5sq�U�����Rm���g�+k	~�����N�� cT��n��wX�'��.���,��vb��kO���]:��ܳU���"��Q���b{{�s|^��&FV�]Wz|fY��ٮ�ٞ��S@��-gSN`��+���}���h��{FQ%>��u��"���:p�䜙�7@2��E[����#��9m�r�ߧ5!��J���V����۬�?�#g�)/#�.ȥр�q���8�Z]~��{5�vTGuN�ynݭ��7�� �^�á/���n���s��|�aE� C39)+��%5A���B��+6�֟�<H��h|Y70c��������r-��ee�G�<�E���g��]�Wxd���`N-�����O�� ���ysؖ/�7i�-���:���g5=/���]�UX�Di��"�DA{>�ߧ�FA��"^,��������1����*Kq�����H$�	6ǝ;*�*���ok쯛����!q	��5�+4���_���
��tI��VxR~6�QF�J��
ݮ�
#H ��M�o'�44���I�וּ��$�L82WݜW\�&�"$]�R�O��Y�� k�Ý�H|!n�hZ |�̖�wHݬ�Ug�фt��d^�x��525�T��i5��i;R'V{��
 ���Iٓ �/q����,��Ҁ�y�@��� �A( �{0�!r鍈�m$,F��!G��D�b忎�q�۫��+��c��*�e����\��?
it^M/4R0_qk��7pq-��v�0=o-�Q�{�>��q�,3��f	�%CX���$���Fqz�J�f�����6�ڲ5����>B߉/CENd|-:Qxm�ǆ����Ҏ�z[ˑI���<�W��J��X�VG��x�횏�r�� �p��6%���(U'r�M���/s��j�`I��赵d��N �QK�3~��\�y��0Q'��[���`�4�;��3},.G�|��G����6.�z!I)]������_��O���4�Kõ��x�rm� ���M�R=?����b���Oq�'%y[}�${��Bu�
�m���j�܄g$?]��`�-����DR���#�� YOc���ڳvn\��£|s��� �,�O��@���E%yѬ
��n]��A�4�v�җ틮�Ǘmi���?7L�LG��Ue�FuV������a�3����F�H�n"_0�o���'�[���*~4�$N�ڽ:��D�Վ�	�E/,S/��ӵe��38�'2�Q�|�~��]�'kb��!������F� �b�Z�ŭq}��t�ɫ[SC:r0��x��h����I��/�l���Z��<\{W�oC������"�㑽��$��-eN��%Մ��=�ɰ�[J>�wZ�b!6���me����EmV��)�H�y�	2�#yָ�FU��Q�˸��5�B��S1h�(�#�m6t)�]�θ�?�Wn��ʥ� �+~�Rj����[�J��N����m&')�����Clo�c���L�����A��Lp�v��m�8��s�&C��غ�܅���1e�/���F����=�dB��c���\��n%�|䣛��q����'�����)y�#�I�{e$2M��w��\�S�a	����DH���B��C����Hb���>O\X�`�LGKt����/���M��%G��h�.!�-�.��Š���`��ԧ�A�]rR��`5	aI|+Ih�O�0�vǻ�jXC��Iȕ�S]��<�
DdA�u��[���D�@a�_�i(/X��
!*VN^N˭j�E�B=b�j�m?%�׾�߯���$n���X��K �}^�������`,����S�?�d��g��j����@�p��)$^��@��;����ٶe.�=e&�f�����h{k���-/>�:����s�>#|y�W�X�����/@	S��k�Ҏ����v��c�)�,�z�'�,J�7��qse��6��\x�@��9��|;�o�ן������d��6��"@s){�)�'�����2W>c0-�+�L��l
��-/��&.�T�����AmWS�3�m͓~$0m�^9��b��?7����5*2?n�<G�ɼ�B�F=SDv��>k����'z���>�Ϧ�(k�X
�=�z}��v��/�����
p�ـm�b����[g�d���wP��LqX�D��X!��2D&,�w�(.�n�f�@Ir3}Ru�� �u��pY{o4l>��"��Cۭ݆r��W�|k��H<�b�wa_��H��o�%+s쏇��.��,ʁŚP�B������^#Ï�V�7��`�E�E�5!m�4�E�s{��D��z��*_V�-'��E���[��[���WE%��nqK�R�:\9�6:�L�n�H�#����{7���=gQ��3$Ã..%TV����}�Ȟ��8�~ǣE�7XU�
�B�ލ�pδ'����f(�T$���-�}0��Ґ�Z}�3=�M�`40��W�1�9}*�J�7Z�NW>?KG]S$\uzj.�3�)�.�>$9�B_�	��	/%;�\��Ի��l+t�;���)0�e���1b�g��vG�a9Aѕ(3��(�]*��y��8t+
J7[Msix�&��*�f�R�OO�ˤ"!`��
�g+\U����o�?t��A�G��;dz�:���1L�zP����;[@�@[��P�%�M,<�Wj,�3��VRC;�1�2���g�������� `��﭅S��ӟ�Ň��U=��6%�����7�v*��&���Z��Cr���/=g���\��~����zԲS��� �l/�|QQ�:-�:���'�fY�c���r)��KҫH�����Ʋ���(�����5Z��%�f�@��J�w~���F.DҔ�
�k��Q����}�, �ӫLWYL�Y�s�&,9ڻ��f�1�^�oFx�n@�ݍ�I|��1��8&�����rt'c�J���!0@�d$��g�f���)_Y	�c�D�+I�z}D8xU��{α?L�a=>R�=;���=q�4O�Т�
�<��Z-���:2�wU�t�#߻�.HE������U7j�	����	G̟Bغ�c�����P�I�i�?����4�1}��)~�Q�4dN�)���:�WP�p�m@�ʘֽ��ġ8��o�� M =1G��t���K�1�6F*�rT�{����S�R�z� mj�޵�b�
��ʅJ�ا�f�&�s��~&V&�fN0V˟߄���F5�*Ɩެ�J]8��ɧ��F$4s6�b���x�TAa���6Ĝ ���	@[ES�|K�dA�o���j����6%B"�.�E_��;��I&z���G��FΠi̫6���t�4�\&���t������������8�I��*��qȹƎ~�{�Č'�ǹ{�T���r��b�b���F!��u/������/LG��#�1�I
�D��6�Q�! c��>5'!_G�a�(�3Aȓ:;�ob'\zy�����:XEZW#�m`t�� &)�p��cH�;.U$�䆳7U����99U*C����K�rv݊�U㘖h�m rbc�ƪ����b5nr�z��0�E6NF�9���6���	RSH@�d���Gc���d�dk\� {c3�f��%��U?�w��W<�| ���Aq����0���~h-�%�lPh3���/���<�P���h6�+����|���r?ntC��#�D&G�x�����W�%�����v�f%�d֬���0r�~��õ�!��~�n�*ۮ�W�����B<8�XvK�e�ݵEY"r64C1�;�{�}u>)�9Of�k,�	��s"{��3�"RP�ϖNUv�~�]o=iJ��}4m.F�Pwtf7B8e���#�5!��٢@ �~���?�,��>���Y9�f�����r�U��>��p3�3(�������֞�.`�6��,tRe�Z��(�.S���q>�z��>z�����C��7���lk �t�xŹ���>V+�5�8��Tj��JR'���]���9���݄��/j�O���h2�{�A0�36�8�1�+�� �zo���L�X1�	���=;���>�J.b=jzi��p�����~��9�z�Ki���[_�m�h�c�<r��&t��@7��u9�"���s����9Ύ���.�n���L��I��ű�re�Գ�ڱ���Eգ$B��r/h�����?��F�O��M���R|�K�vBQ�t�@��B���P~!���3�
t����2�!�Y`Ė�$�C`'[�C&+J5��%�'�?EO��u,�g
����"��F�Y��A���$���A��h�4�쬠�\��/� ��8l��H@���OIqU��j�*M�]f�AbzF��ǱY�ތ��{�e�Msg�#�O����ܞV�*�s�%�ګ�_@b��{J��¬�/{��f�#�`�N^�sG��K���������h�M�'��s�P�����{ �}@����éuķ2��^��
�z�A�3-�uQ����H�zr�V�ڏ'��V�+,����%:h�B�/�}�V��0��l++|8͎y�N�~��3�_�N�hf�f�?uK�nd���ъ�Ξ���)�@%v>�yR���X�6t��:���]T���E�i�m��۳ �*�0�ͻ��.�?)���F�@*J&$m��X=yB��;_JC�4.B��~�	U�˛u��(�Y������Y�{?��r��RJ�h��(m89r1��e�SN����'C���U�n��@*q}C< ���l��������k��M�P�����O�Z�{2��B���<x��m��6�s&6�B�?Y](]�ޡ��w�K�������7��kΪ�v��w0������U�V��C�
c��/^����!��M4�6����\|�5d�.N����0��ڢZoI�]�y!�/m?�萋�C��������-�ÅpW	t����ܐ4Rp�����6��w7�(������y�!y����1���|*" �`w�4�tRH�� |�3DUl��
I�=�+��]�8p�� �OG��9-�۷G���1RI� �	��s���-�+{�[b�gΙ흑#�X�b��Z����7Vph�@�x�F��<��h�83*	��Le6pF8Ao͸!U���ջ�����N�+q�9��@~�Yx�r�:Źs�D�������*��k\�	*g$Dv��>q�:��:�m�w�UV�c��B��a$����[b�Ҏ1�)�F'�w���B�hM���/>���(�	��t�0j�V�b� �e�'�ܾpK���d@�R�HIc2�Tj[��燵���m�>%f�wy��\#����v�;����S�W�ьdӛ��-m��.�/;2B��*��aV�M�8�|���ü�������1Evy�Rr�\����e�r�\.��
��-��QD��)�3L@������1w?��*�w�8�(�r�:A�+L[$]fSvV���j9�1(���L����^Q��R�sZl.٫����$��^dVr�7Ս9�Lb�fV���Զ-�r�g�"�z
����h{V5 ��<3�o��4�G0\9)CY�aEQ2m�<]lHa6|�oL�S��ـ �/>0�úi�?>�-c=�m�i�/��lF�3��@.���~�d?~����&��Z��;�D��k�QT��6,�8Kv��u >;�G��ѡd�+Q�,D� p�[��Ԥ{�Z��3P��٬�׾:۪��ڠ�E+7�L���x�WqP+[T�r��%��]��m�����\0=q┡���gcЦ	��%�(�D���hf���ӿJp������@k�o[��Q�V�� ������<�M�^�5�y"̾���^�I=�������#kBJ ������Q"kװ�M��mƚ$"v���7;+������U/J��v�6]��x:<��'�=Ko��$����cї����Wm]�)!�г�o;!/��5��|� u��*���y��	j}�A�{٫N���� 6:
Nj�L�����{�=4P��|����N �Wx�ee��Ȳ��)��ο�&��Ӝ��V��V]p2��О1:������� �k���s�?�&��#"I�v��/1��KM�- �Vf�w�Q6�g�f��]�/�9���kE��uT�}�3�X�`��u��(�>�-mˍp�\Bi�ylt�n4��k���fh2�aJ(/�Y�p����}g٫��ԙq�O*�+'��|��S9�����;�"<%�\z%����k�m�Pm��!���|�G����x!���qs��㿝\�Ύ�hO��ۭ��q:�qُq��+0��?�+A<Nr
����E����r��������0\�
'�g�͜ �][���9���er�����~*A�����	�U��2�O�p`P��7-��11$"��
�F3ԁ1�,z��əjҧ�u?)/���a��d+4��j�x������!�Z�3.��W�P+�O��Nh�R{X��e�[�F0�=��Vg���f����d�S���Âch^������/��ۏ�0,+q�4Y�k���*�>��[DP_�T#o5���� j�֘�;��)��wƿ
;=R17K9#����Jʈ��WiJ�2+��'öp��T���j��G}6�
}�K�����臿�M�bI����l���-lc���6�H�Q�C'���T"�@�(Ő6���װ���wh��'Ys�̣����T��$��j/.8e0�G�����d%�w%�9\��ho@�Q2��T&�A)!�q��C�A4��%�%�hټקG䬬��Z��qiY��� ]�	gĕ&���o.��=�0������Zg��`M���S�Վ����C������@�āL�^þڌc�o4)87SJ������у����b�y���y��R��;z��w����~���T��^YN�䅇�8G��-M8�i֑\+�zN�4{,@�lp�����Q�}fN���0J,[�����85!��>�4����
�(<y'��*BO��?}�ٿ?+Fl����x~c���4�ս�a���-��U��یiU\L���M($�<0܁;�����e(��S�S��&M/� ܇3�|�E�j���[C�	%B�\wx���ZUE({
xRs}��e��X)h��F�^A^%	c�c���DfJ�[�z��v�m. �GYX�~LX��&������	ԃ�H'�ÙkO��G�'\�<V6% �&���������\117��� %��y	��:�J�
 �z���d�����E�-h���
��e��l8��Zķ����g��T���q7�U;�w�Ia����0��V���qD��w8��y�{/��Tfdzn�joi�[�	��矯N_i�ݤ�T���-�^��}�ʭ�˝g��l��l�XU� ��;%���>��R�!p�S�u�Ĝfv	�1����d�ps��'����*z�nx�YV��ͨP��3�e���m� vЪ0��W�~ev�c�Q�%i��<U����G�v�4}��%[�)��IL���	��x����p��j	��_�����?2F bُ@�'�0**�����#)y���h��Wx8b��޽�زIe�Ra�'	J(ڙ�-�ny:���qO��!��U#i���L�t�AlhP���r�?�j��@��b��ʉ���#��~)
���Z������ ���  ���5j��N4З�f��J�*0��pHoW�E/?��s5D��RN�������K�B�/m�1�Z�Dbq���Vs, .��'D�����8K����OY-f*M�0],74�ֳ
ca���gd?��~L�
F�-=��z�A��7���dq�e~h���Y�M
��!P�d�]��BYI&��
O������- Q'�C(,�5��\��*5�u�4��Y{��|9�R�Q��k�l��^/!1_�}]���QxJܻ���P>z��}��i�"�Û0)Z�}�n���34�.#��&E���f�ኯ� ����m��Ca��h9CF�3(c��!K8���}i=D�lA_�`~������HRoކ\��*R��'�X��X�-]�p;�K+v�s�*T��d���b�g��S�r�rw&�9�O�}��|�Ȑ�^D���b�+���(E��߂�dt��^rf��:��LH��ϔ#�q_����N�b��~�m�Y�j��O�"��~8��j�@.A">ЅK�E��bš �!�\���Q�&����#J]�+����@���O�k�/����r�T%�'�_��)$t,b*�����d�+Z��u�չ����+3\����ș>�i.���Lr *���Ȉ)Le�;�kFmoR��cf^^�@Cu4�V���d���6]�j��d^��mN�ʐ��!�c�d{P\��Ym9D�
lbE�.d#Plt~#.�d�\����O�&��"��ʃQ��i��D+��[|�_j�D{ӷ�å�̪�G�I���[�ԍ��~iVF���D��d����\��&d1Q��~�;���I���"b.���FP��+��6QZ�6_��6�N;��TSQ��jj��>���6�"q��Ž�&ŧ �����MR*X
��:���;Q����c �A���kI�A��U�y&6��M|d�y�>@��7|S��ӻ�*d�P�bN����"�>*���Ԫ�<�5���0L4�yvGf�{��Ζ�
�׊I/Rf�m�B�3g��*�"�Uk�O�+�C�����_�5�=�R\\�O����D�i�i0�#�k����y��OB `����9p�ح>��������,����_��Ӳ�ݕwp�<��Ę�g��5���� ��|��F��~��ޞ�;�:��y�a~<MC'�7:J��ʺT\�
�|)�u�
*^n����N:�Ԁ��H��ֺ�7�h�K-��<m����p�0z��'��~�$Y���X��[X�Tu�U���ӡ��UJ`�/xW��F5>�?deDf�d����D8��W�]���xN�@�8?|Cw9Q#�@�`����IڱM�ƚ6,e�(�h�t�vo#M��f�MR������pd4P����rɷ�Ya�8^�Z(��L��?T���3)����T2
.�r૮����Q棂���$���D&�u[`C`eO뀈m(g��4���Lpݺ�F�M����i���]4�/�i��&x�u(���br>ͥ#�Vy
pr똽;�^D^Н:n�����oVJ�U�mnz�h%���B�t�kWwT[��_�=B�G��cS�/�����w$"�z��pWʀ�r"B,����c>��^��c�_/d��d"\����#P�B쟐������icC�ᕆ\�,}&� ��X�!��¾̣3��#A� Ј3��W����"���ك��wy%����0Chs2r��<^�wHo-Vn9�`>gz�����$K��ϕ�#�:�6����!E�_��ƙ�&<�	w1�$V<]�Ԩ�K���v�F�|WɹC��E���Y��(z�.
f*6")s�;|�o����ڏZ&��.�x0��TJ�G��na���g��:&�t����Fq$T��oT��v���� ������c�HwH$@,�eˊ�7��ﺪ[Y� ��R�s�(��QP��]�U�����}/g&�p����]�-�~��N&=�)����:4<�B�������x5V36����̈́�i@�o�خV�z~nG�{�R�b(F4�d&��2�k"���
�TL���UK61�ϻ-�4��Z���8}�S�ӟ�{����5����֥!�E{	�ٝ�@)��^^�%���/�=�������x.�O�f|q��Kє�̘)Fw=P�ƴ��������Z[�l�p�E��L%���MX��r��z�j̔�ߠz��ev�[�2��;��$s-5�S�R24�+�63�wV�$���%��ZG
p�#�_��L�h��>[1GۣɍIb"�0�.�w�$F��K��'ӈ�R���A�8�l����;��S���Jj�L+��'��r,�fXm��ŉ�C�/no�6�3M�ky^��k��: ��y�4b��2Tj����{��Bn �����_+z`5��OD��'E�2z��ϛK)9���PTS�\rT��gpQ��m�>#2�hԐ�Iz�9�����z-'�6X���{M6  2bN��I8�#�Jk_��P'������VH���w��-B�A`M�DI��i��&�)FB�F��5���o�l r��0�'M��j���rѝ�獩س���s%m[m��y��i?�$L�F��D����M���cK�Na��RM�̙���%�K:��v��Vj��~AvL����/V��/���T!���	͹u����Iׇr:�ad|J��l�,2 ���O�_#Ay $T�I!� 2q�НHj�6H#���d�4���cm-�e����3�1_0�t~��E�S�T����F�R���M5�Ї���@)��.�O�v�']�7��������I�`bك<�M�Խ.\���|�|�^����_(���U���1��S��]�_�Ò�2�D�CZqJ��Ǫ�� ��q���n�e��Vq��zu�ʭ:ִ'��^Yq���K�+;�zb����?�j� ��R��e��<"�$K��(<��Ë?��8�:�>8�3L��O{8�O�W��<Jb����(7c�;��㙟���z�`V���	^����T�mi.������_�?��T�[�lp��~��ܴڏH:f�o��"�)˗�-��������ɸ<�'L����ٸ�U��Ԗ:�C�/6q���2�hC�������<yS�� �9l�)���v�(���'Q�N����nL�6Y����;�j V�0���+_k�74�ɣ�;�uCHb/�u;j��'�t�铞����,��aB�%v����|V��] �uhh��^T�"�/�z.�3������a�Z������.���qIND��sV�W�]�Gy��;6d'¯v�F��a	0��h��>�f{����� ��1<��>�R.��Yf��)�A�늬��Dǿ�!�tI��8A�8k�cٸg��n�y���?`k��lE�Յ��H��^o�{-Y�����z��
7rj	��|�D�@h�; ���3VAI�r��N�h�]��"�J*Z�(f	���bc�<< 6c��ͳr��x�7&d��0a�"��h<�ڞ��/� ` ����
�" �L��[��v�e�FS�/��73]��i��b�g(_�m:�hVȇ��#�C_?{�����7o�az��ȧ	�No�l��+�'��e�E-!'5`���߽��t3��q|9>�mM����a������t=���؍J��WA�:�^��LBLpnF/��TW$(���G|7(n��N�(��<�
Q�]�&̴e�7z�Lr�����)��i`e�)QIZ̨� ��;�zo�[ҳ�����*SY��NU���P�[F�=��(!1�}�'��2i��a�oRt��R�4�l���zJgzD�E�g�7�����6�$$���E��C*��+P�4��FC��T+�K����Z7R�U��(a��-Awl*"�j쓾�w�<��D��2$���8�4'A}��́3�L�"�������.�/4o|t��}�T�6�{��sN�nv��KW�U�Z�Y-W0��%8��=�ڛ�ĖR�X����g/P؛�Dy3L��QAV
pYcא�q���s�}JԄg3\f���/6��c���_�Ht��V�����N���;���@z�3i��]� �i/B�%Sz\d���7~����;�������%�gnF�Y�9L�Y�tT�Iu�Q��j b���x�5;�
�li
���� �p�ƪG�_R�.ܠ �84Q�j�K��fgg��?F$�ၞ��){&QP�f�r~�TȖa/��=���F|��|��(�a��d���0-\��zg�j�J�3V���)}���sJ��>���C�㄂e���.�t�v/�Y�7�J5yo�9�RA4�Ľ�Ot����~�Ԩ7D��(|H󁔩�)��
�B\,O��^���%̳�N����ؤ�s(d��ثC5n�Rx��}��\l��y�CX�2*y�ެ�ڌ2�)�T���)O���}p�f#vW砨�@�g��"���Q� �g���7���P�7Lx/u�h�
�F�d�ǫh��R=JC��^�sĨ~B���ϕ1�"��a>����=�\M׽j4a���׊�*��V�ߵ�1��m�+�k��q���cEH�h�r%��7P7l���"�/�:Q�ٯ��$�!9��bQ=��T�L�����`���Q�����Q�����>aJ��U�N�"�(-~��!��pq1���剚�4�;�����t��I���@�eB3!�L;�+f�?|D=�����Z�>�c���|6����Y����E_�G��F[�&�(����$����(��t�!��pnx�.x���^���6�?��kd�
n_�����*����4�{Xi�^H%mɔIl)Dّ�(�4O��0*�z�h9�~�P�A@[E�̂�"cWY���J���o�_کo!��Xh�\ކ�G�f�=���iGl;��&�r��1�k�M�٢��;�N��b��Pr�)%�Ɗ]�N.Hh��L�V�N ���dK�&�;��!��G�1v�y9���	-���x�H*��l`|:�9%Ͱ��(*�ΔFꖌ��&��t�Q�8����=����,XN�oV9=�����Y(x�s�*��z�qu���`��j�X�h�|�Ic�",=q�W�8���]�d�Ǩ�yА����=�Rܴ|%�ntz�O*�
MҶ������9h��}G�Ia��z����J����x�ϥ�b�َ)�ݡMD�[m��L�w����=դ���h�a@�I�}�{��(��{F��^џ����3��;S��:bN2�V!Q���{��N���˪W�o�CN�/a��I�k�cDƜ��uu�D4(|n��u{}q>��)��!�Qzu]�#Y��p�w���ae�{�P�8�Sf0�U��6(N64��Sp�*o�D7��Hb\���En��aE[p�ߔ�dލ뽓 nʇb���}��0����L���zt��dh�>{F��m^��ն$Uz�F�3]^���\0�h�*����an�d����P.��%�DGb����=�^� v[��9<^�="��P�����G�^�g�������ɖ��X�C�f���_z'|�O�e��iC�1U�V����(cg�wWo��,����W�{+Ƀ�kX�6j��MÖ�@�u�
C�+ �h�zz?�
&�e5�G*��Aa$�G>���6-0�젬D�~#�
�8�Ѓ�H$������1�G���K�m��:� Z�K�\�xl������T�<���:�UN.�����������A�#�2o��u�r��+�$���
�1+�-��(�5��&h���]�h�|Mi���.�ܐ�A���}��>2�ꖺ��[��%��*P��}Y����$�� �.2P���ޟ������q��n*x4�5�럠yn�}�d�[Y�gB�=~���媾d�i�_��X6^�2�q�y�1;6-�إ*��Se�����+	5D�č/�����R��&�R�]�U�X�`&��[��<wy�)�w�tZ.�.yq#W��u��* K-��}��\�~Nm��,�`�	&1�8/�^l[��!���\�9(>lb�З��-��,�����Z����|*����[S,�d���c����P�pw���08�C��ˠ�y�M�v������L~7��~4X��Ki�2 �Wk�`����e�- x:�>I2��ԡ�+�p;�4�]vZo%��5��<��8�Y�%%��7z�'�}@�q�P&�:�AK�&*�K�A�n-��o�g���r�G/GC\�Y�ny�ը0 /��ջ:����|,N���c�KH	i�0�fT��`��̘;����UW�A[\c�E��-��0:Va�h��Ҥ�N܅���	]>��Z_Sk<��p��;h�q�b|%U����(�_���i�����	b�,��+@ǪlK�	�Ī.����"5���en<E(|O��+�z��B��`��Ʃ >�W�1���m�"u�<\\TNW�QY�P:���c�g�!��?��ŸϤ��6*�*�7����p2@~>!��	@��ݸ�;s��v��zUH��c�.�mf�3ť�E�m����5�Q��[����e�ގ��f�9|H���}o6���N�.�+J�6^<j�X����Sx�x3$�����ʹEcw'/�Q�g�\^�f����t<WVS���~:t��V���'�W��%������K8��m�e	�*���G�އZ�I��=���6s#��3L1�k��k>O�l��@\(�H ���_]	U!I:����܃�k3����Dv��s��G��{Vv�2#��1�?O3b�<�6/j���x�o��y��O|*��KL?8I{�1|�]�~Gi����뙢u���*��b���\GA*�%s_��>\�݃�7e��4�2���h��'ԧV�ظbSw��s�:��l�4��B�bݾ�V>���W\��ZءBe�?�����!��K��YO�g_b��r��wv�P75a^�)���_�(	
pz�>��4��y�,K!Fu����@[�0��E��Ą=��� ̀s��X�ٞ��PBߟ}�\̔�V�������/4{W��~���v�Uz���h5·��,��}P�׾�5mD(G��PWa����9uO\�]���]f�_Xq�蜊�Zd���l�t�8~D�����k�#3ƌ�jep(�Xo/�v~�tF�l��_]5O�Vt���"��_�^��8�Yiݛ���F���Eџ���%�t��d�D`���
%i%[8�x��T��V�ü�Y�b�y��#<�=���H��Iw�P�r��$nz�2����m��9�{��.��#s%pq�m�JʶC���쨈ޗ7�eJ���\hE.!��_�;�W�Ĺ�`p��(|�
}M�gXT�¾r�����A�1_C��B�۷��<8�Cꋩ�^�8RF�}���k� �|A�?=���f�T_�� j��G;b1� �������Kr����B�-�u�$$ǜ��m���/UG��XT�O��lՎ!�H���x+��q�d`�*��#���	YPS�j7�Zj�@�����KT�ʜ<u_���'�0g��D���93.��^Q�)O����K�ۛ� ��9���c;MA<�Ks[g	�L�b_�K1�U�J�w�p�_��bSn|��W��N��;�Hx��A�R�(%�ND������d���h�!.�1!�=tv���#�.�8L_��
���m*���{{�+Ã�M7��R�J��7js����݃P�oEY��a�����I�����Z���D-YXZ"��E���T^�r�Y���9�kt���A)ʹ����aW��	�����+�IK�P�L�O\��V����)?�av�Ebꩠ3)7u;�Q
Р�}�:�1�+�/�6

D��v:s�&S-su�O��A��`Xv_�8&��r�b�){e�6����{_ȐgM�����kr$Ȫ���E \j���`���C���Zk�p��?~Ԧ��i_`�<W��"��ǀ��.y�2VgM~&�F�q��?�ߩ���M��T�mx��'-��#�IE��0Z�YrEY-�F�fN�9�{|���jw��=륫X�i��1.Ʈ��Z[��P�����ٟ>�[��`���P.΍MVw��@�4��8_.�ͫ�Y��)�DC�E<l�L*J1Q^��x�}���+��<��_��B�OJ�:��9��i�Ŵ�z䗰��n*��)������T��6�IP�=`G«W��H��1��<-�#�R��R`�$�[lgOn4�ko0��g��:oo��ʻ��1��6UB/�{�4Q���c6s,�#"����ʏ#&����	�3��u�W�d!5�s��z�z����#���8��^E�B)a�<_%�S�2����6��Z�ec=�]n/�#-~�k˵*�9,ϟ �����}��Bes]�G����
3�2���ߟż�;՝�x+2�i �9U�&*�����֢���{���6������)j:7��]� �0��0o(:pP���À���Ǎ���A��9$����(K��]�}x/p��[)�c��O�a��ɓ�i�Ƶ���fJ�C��B tuB	`��![��[�BH��*QK��s�k�&#\��@5��P�	�DM4ϳtT����
E#~�}�a�M@�����6�x7+�uRFƏ��+M��I�e��蕃���&s�n�O��]:^�F���۪�o���cKH�S[^�O�^&�{$���<ȅ�D�1E�&5rQӞ��m�(
p#��]Z���V��#O)i����=��g���'S�/Z����g�~T��D��w2W?�v�z`��TP)w��?m�ݥ�u�M^9ؼ]�.ԯ����{+q!�c����緊p�j�E��-��K`
���e���y���U�����B�u��a�k_�ڜoHd��M5�|�cr��8G��'[VTF���|s�:�ű��6΃�ݩ�/c^v�����m6Ī=��[�y|*��^"р�'FmW�qBH�DPFz2x�o�y��&��� ��;���Ԍ�b�qSu�3�`�êl����_��'@���D�D�:�i������/�1�0�ځ����Q��̴����:�Q}��Q��9j<\�@N���_
kY\g(Q�KV*	P'X��W�\L�����`x$�<����Մ���nrVɅ?
&M���m燎��)�8G��	������	��l��5(2�C���5�Š�C� TƩo;q۩ֽF�Q�e)���붩��Eu��|����lӱ�C�;�G]a���H@��&)�琝���ӔK��������f� �W��}��pF��,R=�!�}�cY�nKK�7�� ˳W� ��G�2�f7A`E�yV�Ҭ� 0�A'�䉬l��@��I�h
����o�	C��sDO8]f��y)ܺ���A1	���A��{,.W:Y��+rVQ	z5�����a\9vK:���*���:���/,�Ni�]BuS^<�0-����s�o��mw'x:@R�>�j&%�Vp�5�\���~L�2=1%N��'�Nl.�yA��S_����ps��o@�����Pz4��s�?���?co~Vg��Vu\w_o�b����Ef*2_��g�a ���Hy<��%G������[a�A�\�iQ11��zV�4���FR��Sҏ-j��cl�%��_c��u�����A�| \N��ACSm��	�SrB�=�Q��)߫k��d��?����c���3��Z�ޛ9��Vd�����b˲�ɅMG"��������c����A���%�!�iw�1n���ӣĺP�e_��]�q���\e����o���s�������Zn���Tke�����%����Se�c��v�X��k�[�I69��a�{,5�5HRgκ*�zt�e��DJy�]K���c�ҿ
z���J�dU�����~4?X��{�`�OVOU�����Xht.FOtXG��g��j���'���T�B|�W��e�9�L���z�o�x�ˢQW�Q2�� 9^0�4�ou�r�v70Mh.Z�����.��Ͳ�h����2��r$�a�)�SU�<���+cYuב�9QQ�$R2;�7�%s�7a161�UweE�]׀y)�[]��+k�'��]�R�I4�>t�� 
M |��es�U{U��X�1o��#�8�*�׺O�7��j��إ�a��*�I��F$�,A�"{��]C Պ��
���7v��N%��U �~�����8L7\�<��v^#d]R�q�=`6�ẻ�LWPjЬPl�(.͡ ��,��*�X���5�b�>AX�d�5�d�I�w(j1�o�nUj�l�b�%��H?��6�b�w���#�ZJGve�J�sȘ,� �vm�s���Wƍ'�\�q��ͿTsT�R���o�]�]�y]���a�]2�h$&F�q���hI<ďՎ0gH6/d���T���A��T��a��J��8�4ϋ������ō�j|�˛=�R��yW��+Q9��:�<!`(T��u;F�?�'���5����2�r�r~ۇf�.��^�9+*�G»��6S�	�L�k��
%jm�>��D��X��S2���Z�<y��^�;�*�x����K��Q�n����=����ٌ>/�X�䁷COP "��6��PY�����z��'�:/��
������Y6E6�S���?{H�pDǑ�>k���{8��:�)*f[����d��r/�4= g  ` $�oDpn�	m�[�������n%Ջ�f�>�ysh���$m֫��w�E*b�t��r�v&lO�"VL�t�{3��v�#P�s�`mO��c*.�+�����N� /��ʝ�e&����l-�g܈�[ej��c�[�<-�7�Ht)Fk����8���� ]7o����.S�*�Ƃ�=�IF����/7a�������z�Ɇ��~f�f���o6D�A��_���B��a�p/�}O��w���nZ����0�[��BbL;'�2��o������i�*=�S�"���z�'83�B�6~b5.߀T�8䇛;U��!L�@�֏�+�h�#w\��o��0(�{�zB	�0WI9{����0i.�pٔ��%ő~��!Cv�ȳ��C�:�0W�h�F4	g�Zp-wW�Wa�a`[�dX�@H�J2J�� (D�~����)]��(ޅN�DB�� �E	6�y���g�+0@��R��=" Tg�]����=��Ê�v����`4�H91偈+06���P��{}�F��]��a�V6;{����=��5G~<�7���X�f��1�Aw<�N%��K�()��:/���C��w�1��E;�g��8�[O�e`�+��M��nG ê`n5Ԑ�	�-O��F��:�r����Fҁ�����R����:y*�R0w���DfsL���h������W �oǞc�S�[�e�Ζ��q��t
�8���5��hǥR����R5�E��2�il0=,7�`6�t�Ǝ���뛧�"�\䩀�HC�����Ply�!a�Ǩ� ���"�/ປ�4N�4l�/�Ӕ���e�w";'/mTi�[�'̸���8�	�y�s�s��x`��3�r�^%�:�;C��x�W{�ޒ��t� ����ш�x)Ԭ��m�S����i)K���HtF����Լ�}�Y�� �3ԇk��9��e-�'K ��x�F1�\(�E{PV��2��r����б��;�x�]��{��sK��	o�O� ���v���?��9E�A�4�&�J/귧umJcĬI������Gd\1���A� 	3xb>,�����j�oM`�E�*�@&��A�a��m�Yu��V	��8��!/�,�P������i�i�^����t�3�R�ֹ<��%�l���lWp�Ɲ;��1���$�YR?�=X���%�{�%�![���Ѩ�A+^
��<5k�������Gru��Ϭ�2Z�P�u�Zcﶼ��!l,ν�H�^vH� bIE��-7�ՙ�"�,NH����G_�>@�8�ȩ-5+ ��[�e��{@����\��9�L��t��o�6L6�p0�h��Pmf�s����Z#a�_KI��3�a��jN��bĈc?��{WΑt� ֳ)�1dx��~	���gB�,�X8<�g:R���-�ɩ��I�G�T
}S�}GէdS���B�2Y��C}��7{=w����V-�(� d�D�EZ�D�^���6�����S�0���Y�c�F���ݷ��&��Õ����횊������lGG1hXX����&j�)$m$3�_}�3p����})5�"�����bnB�M��\o��,��,�=��_�Ф�W�y�O�;��D�ʬU��M�a|Ҡ�����
9f�{=����T��i4��̣���jWp�whh�%����6?\�[ͩt�A9X�I��E(P�qK��w�J�/�γ�T��1�Ӵr����]^�>���k'^�g����b�rn�;l�^l1�<�f��Q�> uoeE�`N�����R� �r߲�w�P�]~ x�T�<Q�˙�y��j,]䐿��%��[�>�������
�T�l����xEe˄�1��><��qb�����~Xq3�d���˜����#.����!�4%���2c՚��5�j��Do�Z�):뚷����0*��8=�j�*s$��J "��+B�LnV����O3[�P��ܬ[!^?&�N�?@��U��ɿ�e�����O_Lxce����[M��IX�a�
Z�2N����$��ZE~�ԲC��J쟗��i�i��~���^��Fm�y�+��]�8Z��y��죏�2�{��~Ȍ����;��5z?���^zf�=i�D7db�V﹍Y�A!y.���e�$�u�J$S�e��,��7��3��� ���@�Y��2?yr
��b\�\|5��|2Zdl�{/F�B<Q(�_~/tj1�nb(FH�$�K`p��9���Ƙ�q(�'wJ��`�5d۟5�e�?�C�a��--?!$2���E��(�m���v�uKq��@p��!�L�x�sM����0��/p3�_��m�����Q���������>��RRuO�
q�>�r���!��9�D��	z�-���{��ѽf��\G��.hX��^1G~���\����*�_#jN�y�ȶ6��UB��Q�}���<1�� ��T�>����uN�h�%�d���1�7�tqe �1�]�nR���l��ԡ)��u��D�ӟy}	��*�PRy9�<����..Ey;���(�_�"<�M �w���e���@bI0I����I������`�hSw�F���v��s�k��L{V3WǱ�l^Y+�J�p���Lpm��ﻰ�q�.[�eaN�ţ��H��O����?����|���,R6Xϣ9Yd�Ң�t��8�i�<Q��lg��)l��!h�K~�2�_�U .�yJ�����Q�O�u���h�n_�;.�,��A��,�3�-H�6�Ц��_��<Օ��o������K�n�z��j��T�s�o�1��o�Ƕ邲#&�[]��F>�U�G
{B����|�t�йL6�`���Y���1�jG����!�&� �a�y��?�G��,�tA�� ��Ȅ�7\d����_@=x�/�K�'�f�͸eb:jC�����7����H:�����	��֑�ΪY� �˂/��2�b�!��e�3[�Q��ԁ��G�j�b��Uf�K���s�'o�ʻf0���E^�0L �BC���y����
��A?�%��|���W1��H��i^�]1.Ew��R�A���gk04M"~\W�����ΧD�q���On��*	�}'P�b��˜C�?AR���`��ʖ��gY���ԫg�es4R�vd��w�0���H��z���n*�N&J�ݯ��[M��a��;⫌[أ�+��Zv��߆�, �/'F7(+l\��5��k�d�Y��ʸ-��l���ވǮ?�r�����b$����!�F�t�8��z�Ϊ��=Q d}�i؇�=�߯t�F`�p�@I�T���cBs�Jg��#��@e �ǸD��vz��nY�#޽�"1���޴?�P�Q����2�����
bw�>�-H�l�����f�O}Wឩ.�ФŽP'<�u,Lc'���}g.����F/��f6!Iţ��K�����H ���4�b�
b��Y�� ?�ұ��<Ť�L#tAL�����{hK���/�6�6�UŔA�|%�w��Ɛ�Y�ȷq2�$q���)-�s__8��V�m�6�3��Ӣe��?�n��_u�nH�TGv������`��v׀Z�RVp�wJ�d;�����S?\�g�A���3��1����h<D��UL�M���R"�,Zv��a��Q��Gn	U��=Q}���D�V���0UE:��1�VX"�EU�^{���Q�~�i��ͳ�����a���A�w%��!�� H�;Z��)lF|��/P	\��D�@ի��/Z��|�;������5�����1C�"��%�"c"\#	i 0��)9@��W�՝��"ޙ��gD��/�����=^�1H/V�dTi�[^k�]���v�.-X����˦�zќqT:Jx����?Uc=�	@Zͱ�U���@�[Q���y��UEu�_�_>C�K˻�C�_Q��)�[�e�s��l�;8�G�u,�`K�wN���T�0�N���)��Ri��ہ�8��n��y�i�������H!b����u7(��k�D�W�<��e��B�����I�!{sy���ɹ�|�aq�b{��i����2�ߴ���Uh�a��nI��j'�Ց��9������ fFb�P$o(6��ap��G�PwE�*�8��@�1��/��RX�!XT���l�,�AAQ�WKb��k�U�"Q��3'ɞ*e�����࿰HR����!}�G�Q܂�1|룫R-���7��bҺ���+��cSz;V�А���*�����tl�	�yY@�����DZ�-[;)�5#3�.���9���rd!<&����H7�a���6�����c��-��Iy��#2&�_�H��_�vS$���$ӈ�������@7�mS�<%X���s��Y|0�}���~��|����ŧ}W�"�h������3�=��h?���K\5C��;�3����9����5�gZ���	�|���9�O�ƺ�@+D\��r�d�v
H3j��7���ҷ�����p�E��U�'�;r��e�\I��߲�C�D��6�����ה换���R_0���e69cg*x���!4�k����M�}� Q=\D	8#~� �G�r��U"�����N �WEO������V��ZV�# ?l^�6���������15�X\~�K��D�I->��4C,�=�����x�v�&��Ԧ�XIX���}�bT���*�G��~'*��������n�AU�ع�VoK�`;��&�M*��X��yɜ"�؅'�>j6%��o���]Q�L��T:��G���a6m%��oV��j4��Ca>�.`����ăpσ�$~F��qp��U0�/q�V�ᕢ9�\}R��0H�{�M��=rJ+¶�(!z`lw�E;��4��5T�X�dy��p��-(������+���� �i�FWiU� �.��
�D�C*�yc#�d���H��ȍ�l.ȅ}f|��V����Y�~U;��Ԕ���&��õh$f�����hn臷�`���B�so[{����z=� 6p�4)�Lq�^K����gM�ܾC��l!�j�V��?vs����%��n⁸xR�ū�?�95��%��7Ǯ��)2��w�̎̕�p�2��N�Y�� z-��+mu0#Z��{�-'L�P5 ���Łb\�7�����]�/u����J�]:��YpLk�Ҧ
��ܶ=0��H���ׂ.@+����w�e�%��"+5�#�vLS͙�侞څ{<f�m�8��+�~��Q{Y�w#��B�kRn��b����0��{����=Z����Z��x�%�V+��J���/9�`v���[�VO�e�#���7&e�z�[�@������3�#TH�y��&�a[R��
��{��M��Z��D����#c�@�Æ9����K�����H#���s3�W�XJڭ1���Z���X*�
�xpN������9��\v��C,뛵�{SbjDrB���q��5̈́e�`ق��d��>�P3�21`H
�t�K��Pg�URA���P��)E<y��uc�.���P�Ң����?��w0Ǝ*����Dbw�o~����j�4��3uXN	�B�tȉ���ߨ��� AD����C< 3'�롶�姢�q*yP�n9A,�|�%�����O8�ɢ|*>�T���Z�{4�B�ˣ��zF;-�P�|C[Cl;^X�����ĺi4��"S����n�YK���kT�qpt��^��ĩbm�-�J��m� ^�����tN/����B;G���j�"@��O0�_��V�T��C�:Y�HE1�i�
�����	+6���V��샽_�d�58���Q��z�J���O-t�ڨ�����R
�ݣ��f���4�vw��P'�r5,����d�PW�V�)I�nP��S����1j���>�����,�4uHQcW��z *PSr�Q�Qm��������f������5K���BH+�k���ɑ�'�/G$����A�D�i�e�ɢDGM
�'X0�~�K���5�v����Hk��Q�D�<�:�/��T�dȀ$=&�"�Z��b�
f�(uu���|����J����j�=��߾I���2�>P� �,���B��>-k&��H�@��'�*����'���i�c����\�#�W���җas~(\�OQ<7Z�A`�
�������X]�Y���G-��l[�_��I6���П���R�P�f��FF|&q��MG$1r���M'��l�IwJY�=�޳M�<nܨ$��8�n�/�͚b�ԍ���Fډ��%ţv��� ����$(މL�?'��}�S�	�֊��J���vu_9�}�I�+��H�}(E��(���e��Zµ5��J�-�o�'v%`�m#�if̲����.$��&���Ҧ��:�Z��W:�8�`�BVaآ�#O��o�)!��4�c�s��<�F�ӣ�@OX"����t�p(�3�Pr��P��c�HZ0-L�B*�w8������� UKH�-/n��W��V#/����;4���9Ag/��= ��F�A�k�Ⰳ�FtV�m�|�M8���H0�F�G��+	�h|�%��5E�������E�1��tl	Tc[�,݆[`g[���?A�@6P�>!&B]o5(��p���Yb$�� Yz��!3��_l�����W����}�i7�Z^z�4�Km����%}h1+ۡ8޴�Fd����z���1��0:����Y$	��?���u#�C�8wIY��YEa�s*c�'ܤ�
���ڲ]���0J�Hr�P5��$�����Z�V\?��ߦQ����
	�D��gō `_�e��˕��z��2g�rஜŢtB�@;םE����"S��"wj�ri[���Q,�����c}/v�ʒk`0�F�~vk����P;���Tm�I��ҍBQE8~�9�'7�C ��j�^x�7�"��ȃ�X+׳/mER�W,�W�(e2Q,������Eܯ(��yq�+�V�L��2^�-eXO�7���TAѸ5y)���g\eYk9��}H�P:&ߑ�<�G��E=��_�@J�	[_ׅ�����
[}�� �
�ٮE\<̄�G �g*��g���i��Դ�%/>� ��������������y ��|�ʏ�L�>x4$�m�������R�X�)��jY�����>��h:[�d���T\�Lk_�Ȇ��
�S߃�@�"˗���.|V� ���u��a�9Q 7�@j�=���f�����#=e M���v���e������&C��K�Q����ݶx��Q~D�*�ޅ�O���*��!r��I������C&�U��xΔV�
h���܅Xe��W)����؞gM��YȜ��2S}�<�Q>�}CnϨ	Z�͈ѹ��U�Ꝛ�:��XWq��C呏d=��g��}�&>r��˹�����o�?mHk��}߫���N�d,�r�i#Kq��Ȱ�0Jo�9�Ѩ��4gr�*-SɝE5���	��_�=�cmw��X����-$����'�������&~��Ǚ�ס��R���^��
7�}QJ|F8������7|��i|����������f��'/�JXy-vqȢ0+� ,�<��f�;�m\�ȍ�X�p��|��Nݳ>�7S:86.�/K�f�����	֥�)vd=W�ZfLs�F�,r�,U�.���t�}��T/'x�Z��Z�Da�8D�K�5�y*l�&7����ȗ�%T%J�Og[Ԯh�b����f������	��0�BZ_�P�|���UFT��Yt�u��7�MlM@�{3�$��5@��k'�Y���󸝼�P�����G�<�c����K�������zA��e4��7\��&��ã׬�[8�$��+�����e��C�VJ�y����b2��fH���g_u��;�)Ȋ��?�� �D�_��mz�?�i-1mB�
�K{0l�9�&���Ų�9��q�a��)���E�c����I>,�I�U�R{����jҁ.��o����j�]����Ў��w|,�zM�cUcu(����mh���F��A�1�	QaM3ύcp�yk����H�`�7�3#�"m���e��4��X�l5-.���������&�pB��X��'�E:�&��>5���4�������ԝ6�~��J������.���T�"�Nh���_�P8��RA���^�����Zf6�\�D_-��(�K�?+��p��8@���i8,�:K켇��SˈZ�B��`�
 �)�5�d�.���06���$��X1��5Z7���[3Ō�F��|�
��WF�"a���#m��(�hF�Q�Y:*Ӥn�*�,�����˅yыbqTb��5#�=��r�lK�^��{�(HC�X��X��	;�d	QeZ���C�WK�L�~fw��}��j�&�j��x����^i��+/��w5��^n�f�n�x^�Qd>��orĚ%�C����p��N�l��t�>�NZ�P8 ������H$�V�����|�:X�jEڧ#�SO�O�\��H@fxt�Z����x�EՓ��B�p�v9�%¹ȁ�Vݼ�Rƌ�*3n�g��@���-��ރ/*J�����`L�e��k�h.���:5F!6XRm댵���#^�/p2g���������'��'{�M� ���c8� I��xP�տ�0gɀ��ɝ����g����úf���7b	G���={4��p�^v@w�4��m����)��w��ސD( Yu¸ �!� �dm�I;r�&��c���3�������KE��g�6J�L�6���2F���D3���jh���r��_,����+}��	b8�
�Ƨ�c�?��9���	��Mu�j����gd�y�iGε��>�|h����Dy�}<�6���u��L��?(����~���(��?�yB�2��k���G�Y	o���I\_<��\���V�H��)%[E�vH��u��nR1�4/n��k��Z*�)����ug�p�ע�Ǒv0l�� �e�˒�q2��;�W7��s�:�
��P��Ђ�6�s�%c��W�qqƩ��be��w�iA��"�G��&%Wc���$��ɨ�M�����URKXêE��c�mݨ_p�9���&�����]@�����9|�X���*U
#����j~����xR��r0�`���G;ܺ����&��=˪Z�d�nڞ�3{_�	b�Q�.���N��M�r��*��˨첱�*��dF�O�^J�E" �<�X�tT7<��`�$���Id�j$��8�c���T�u�bRb��,b#�F��B#�	�z:V�Zt��x��Z�U�}ɢ��}՛�Jo�Zd_*v����[8R�o��a�㍂��?W�{��(�V5�|��������>}�|��,���-�YDU<�>�p��t�Z�:���~u,k9	^C�J�Za4�n��%�<hmJ�y8A~:	�BcT��<I^��,�[νS�YaL$�gm<m�V���{]+�g^}�%����C��F�w�x։֓uQ*�"��Js�JY{��^ ?yLc�?�w�"�+q
�P2f�J"O$�ș]��F��8 ����g�Pv�
�1��y�pQLiL���9"��#��<c;�ŧ�"�}��=���1c����J�F	�7e��K���`[iy�*�d�nIg�Z�i�+�ܿ�/D�BDҪ���񖑿UDms���Vu �� �����D-�7Q��H�.k2g�!�O�C;���Hu����bB%Y,zd���H+T����'kG)�m��bo��(�:I$oJ{�0[2�U����J�΂�x$ʕ���-�[G��R�5��9�n�92���.���d��f��`~�����6�Td\|<�_Hb2x�4d�do�ԫ*�4�j P�Xa��W�"�.�fŮ%8�BO#|��be۠�lod]���O �FLR�2�����5�[g#,�%P�6���x�$��A�����S�4�C[�	��3h�)}��I���i��C
*P�E{P_�_vS^�����N��ޱ��4��:��u��U����X��2[���'D��og���ԫ��$�(����`	l� ���_
xK����]í�hlz{t����>�3�l�s'�?B[�����	�<Iv����F��X�!tJW�4n�:�v�U��|��Qe0&ivrY3mrƠ�D�<����HsŁ��Ij���O�:do?�0�b����\�e0���Ǥ�<ah�/�|�B���@T�Um�ԏB,�coX�[���NFX��-]Y#���5��C�M.�!��׿Q��&`C�^��R��ҟ]t������,|V�n�Q͢(��EEqY"4=40�gI��=.�mS�u�A����WL9[|\��᪱Jx�m���	Ҡ6��ހB�	1�
ԕ�-���� �<P��纵�Q��M��c��7��嗼6��Y9г�n��1y�2��q)o�R��.��Qt�v;
Rm�A�:��> ���	��O��6?�%tͯ�,C>�t_�]��m�B%�|���b#Y����Fpܕ֓�R�х��R~�Rjlޛ��Ur[R@9Br���4,�\)��R��Z�zX$As�tG�XeS%��j��ʙ��##��=�u� щn����ɗ���BO��_��u�A�'���b�)tH�>B�:�'i#3�~���o�@zb�ьC{{��5��� �.�um������`���@<B�v�٥�7��&��ʇW�b0䇀g���gb��瀱q���߆�4���c��^9���.?��ҥ;�X?yiSo3:
�z��e����Yh��n�q�B1���TI��;S�Mb�*;,������䭹ܨ��PeU�z�G�An�Un)� G�ˤ�:9��%i	,�%�&�к��J3�����#���qW.&�X����%����D�9'Ix�>�^��X�+L7+��� ��4a��#z�?���p������/p����}��M'qK����t��;-WT�R6���i�KB<�����ꑝ���PWv9�cz�����[��*�H�E��p�		KR͡/*Q>�9��0Y�[p���-D��,1]M�Z�2i��4�f?����ȷ{��?��E��I�?���������*U���@X2��9m�m����Cg�� U�lyP�y໫����1*I�+y�$-E�7+g��%�:i#�s�Y�KH�{7�:*p�Z�mksrp�Qw?e�۲%y��<���c�
9xz�v{~�To' �m��፺'{�K���#i�}A��"	�a���}4g���a�]�!�y�%S�k����d8iwc������=W�<�(��#i?4Px%�E�[K���`'B�=oR*�6E�g��ĽD�s��Va�1�aH���=*��ˀ�-�{�e�{�Ye�D	�3M�3��tsm�őz�,V���1��o�9q��]�i< 
�E� )�{N�}h��xgA�<`S�l~��z�e�,.X@���tO�LI�*�;��Ӧ}���'u�JH����dCr���a�>Ȗ�i=��//��#�%X������FZ/a�����vOTX�CxePGp)i`��*O����.<*~p�!t�(ar.�`?U�.�ӎ~�������c��S�Ra��A�Q$�Hθ�}ol�x��R���W=�_�bo� ��n��/�~! �N�3����1��p	#g;�!�u�7p�h+�b���Y�1�Q|�
ػ$��#����z�.�w844vA�N�}��B
���>
��쏶AX&�ҲmnG�E�qт;��z��`�m�c�I�&���%׀��d��
��ק��f�K�D��Ұ�
ͻ^�u�ke�D��;�^�J#g�ͳXd
�ȭ^����g�Q��6Jy�_t@�8��I���\�r�[$m����89���nP�"�Yϙ' �n'y׳X�	�a�u�o���gpS� ���+�ܱ嚑��b䄗p7��p��)�켺�}*l�0��`�j���j��<	��������f��?LF���L�@����ʙ1튔D)ظ)���)ݝ>2S�y�^~�y�T��C$?�����+�ɣw&��+=�ަz�����e<�x�O)S�(A��Rw@l
Zhy�VȖ+ߺWlP��o�R2qN��)�ӎqʟ���R�U�1��c�[��#J�i�ɕ�O��l9��!���A����&\�f��n-��uFvI�+(:#+��M2郫�%����D���V������4Y�D@2�И�3SC��S�p�ǽ{2����A
F ��TY>�����o�^�Iᒱ>.^.7�#?��n���R ��I¡�t7z�wcX�����1Y�D��U�}��PIu�K����9Y��]=}J�X ���7^������tXGVuPNDH�Z`��\~cԃG�;U�.m0NLf$����B�z���0$I�<Bso���Vgf���	 ��`P�Jg��Jl�C_�7A��gh<�Hޣ�4Q�ѓ�B����X���L���J�7yC�0|�Y�[jFSk�ʖ��',��X�i���E�ڥh��Jih�R\��F��6�.��f>^3�jw�"�F�OV�d7e]�W\�C_wp\u��t �?�y�6��p,������J�î$/��w� �k��~�۲�'�&��-s���l����b�f�������Cs���c�*�|�m�}C���g�x�.��������|[ڦc�6:f��E�7UX)�$i��}ʀ'4^"������[���L��%�v�8������¼�����Hb��9�;/�UV�߭~������f�����[�w�'�-���~���W����-����x6�15��Gen��d�2��k�^�nfev�vu�� �-c�>��8��S��}4z����ȏq)�ΰ��i����.�M��z��k�,fZ�_n��9����I�KX�����n��ƛ���B�dClM��9	�f]����K?���򠯾��a�ݱx@����ŝ�ku2~R��xR��ڱ��jpF��r��p,��b쟙�GE�+�?@��"1��Om�F��Ԏ�m��{�U�%V��#�����~���5yQـ�d�n�K����qk��2Ь�$MWh�����Oc٩�mp~�?�Yڛ�GK���O�ɘ�x�	��6�R{�B�G<1<�=a��::9��E�m�T����c�VT5D��7��f,�
���p�\'A�M�ɯ�Y^�\J�0I�ȩ��;윹�ްk侀,><�ԦL�=,~$��[̈́�����҄]*��\��s�So��	��qIP��P��퐻��V�Z"1��W�CKb�b��^��$������O'��i�pU���H�s@�UddT�ݗ�����Gܰ�g9[��r�������n�I#��k��\e�j1�	r��w�Q��ƹg��+k�����L����Qs¤*)��.9V�a\_��½��E1-����/,{:���^T���hf�<�=&̀���wǖ��X�
�X�@Rn��f9�_}_V��N�A�켺�4�*��W���"�e��lk�+�xK!���I���j�s����YQQ�h�n5M�!�a�C6�e�_�M��;
��ֹ:�9X6�8��H�?��[m�1p[�2��s���&�z��L�Q��D����&����O�y�Z��0��.�`��g��k�i�Iv�m�HM4V�XMXf�>{3均��2B�{D��ϯ�#�غ�\v�P���H0lP�v���{���7�%�eP�,Q�(O�	��f�V���`���5#~���&MҚ7�������B�H�ǎJ�/�f�w���Ŵ��^ x'���t�����i�T�x�������d��p��x�=N���_�gS�?"�<^��o��h�Ya,�bO���'���Ey��KeMU����r���uZo�w�b�Ǟ�Ti@n"�m�9��gR4u�cR�:�F�]
9�r�X��������]H!5��OO�{I/�J,��ܲrA����X�w}�o�"?SF۲�|q����b/\[�=���@dKg���lY��廔����J=��C��`C��LX����Q^�˟>�� jԂ?����|kPX~M�Am�Tq�	H��#+}N��Ո&C�Vms�{��k�$Oݞ�J���\`4���dVR?�ws�%G�	�Ţ�2b�,��՞��.@�����gCI�귷���R�&˔풇�H-a9�ҧ�Έ�+3�1itr�Y~�L
]]��M,�64�Eq��	��7��ߍ��w�MI���.W�_���wo��=�����Q�5�������P(�Y�{�� 0q��f:� &�IMx�^���d����v�!�ĈIةk�0<�������|�G���Jy�Q�-�%*��t�����08Ŗ�_l$u�'�����j�d0��KG�A\�_����,�L�d�Q��L���I 4B�YшO�y������:��g�5u!������'zn�d1��$ݻ��M�k��l�灲���zr�4��,o�o�ݝV�zE�w�)�O0u`��:�h�Z-`х:���lp>��҈���@l!��e�g���P��=�*Z��!&�M�F�&�1j�����yGFG;_�R���D�e�T�$m�5�p��g��M78�-�\'&�g���3�C.y��m�_ �o+:�Mr8�b�ɇ7b���0���sW�ۜ���Xb5D�!�F����ؖTuC
4K��NC�	+T*��E���v�zng�eI�����#����Pw*d�ܜ����q�/��L:rĳt~ß�pO�'�6l���}cp�E�nPu��5xM�Ƥ>�60�u��o�SF$�ܶ��O�� x�?=	�<�����˧��ř���vK&>E����-�PǪn^R�v6��^�s�q����Z�	W�µ�*�z������?a�6�{ތ%w�^弖��V�m-��������n�(� ���'.<�5�L����S�����'j��`N������_��R8��`WS,�[�Z�9����2,�R������G<��{�b��	�n &�lѯ�68�T��J)Jױr�����tq��� r0C\
D�]Ý�:���q�τ�aa�� dhj�Å���Dl(EMQ�?4�,e�����p�?�r�&!1v�Z����H?U��)�n=X�׹���z2��n���f}����@?�n�4>����P��H}6��j���䈒:����ҍ8鴷�QU�?��.%����Ԏɸ\U����{I��[mz��$F�6F������Rt�G�r1��6���fw���8�W���\ z p���]�7NF���x�C�KȤ������
��3(=�<���%�E����B{3 �<��h�U�4Q��Y�U@ ���І�-$����M~��2�V��	*I���	*����5u  ��Yy@��ȗ��ٽ�{TKRTtH�A�q��!p#B�:Y�Xݡ�A�9'�t���
a��Vk�3Q��X��Re��A`͇N"��^� [<�e�!�5B�%�8���0y-y��aD��p�6sC'[����cE��ͱG)v0���7T���W�43��'2@8OSTp�fh�M�u+Op����̙i3�����hpK�	D�x}/����k�X�B��'�,!uv�8
�+����2��괜�0��FvJ�?,��5�jι�?$�C�\�n6�іl �_!���{�LU���������u�rH���	8GKM/x����2(:݃#����Z��J��"�P��Ǆ��%���5C *m���Ώ�?������bD�յ��BQe�=��+Ls9��t�����h𓀜�U�5�w��滂��1K0���$'p~�����ҧo;����5��Ds�-E���8�C�K�f!�=0{�?�Go���xd^��#s����ϧ�y�g�V$!��1!X�+{���yr�����H5�`��^wPl!HGT��4F����α�|њ����f�Y�
IEz#]�RQO�̦'3��oo���/���=U�e O�W���v�W8y��p���O��Iё��هS�I@u� ���m���U�~�m��d�Ή�NL���� OwD�5���o���pK��?���
o�R��nh���-q�<7�h3�Ѝw ����*��(�FRﻰ��.{9�$�EOκdI:��u!��-C(�����F�ٵ�L櫁L�/z?���`���,a�#�8�;	X���ܹ j��r!F
p����&���=a��1�x�p우�c`.##Z�;)c�^=�U���g��~XV��snS#�2��jCNv��pr���Ő��t|�\�nAe�<�T��)�c��*s�-{�7JX:5%$3z��Y^n���sc�q�#��%�;�L����4_t}~fLܴ+&�l�W��6�J�6B!ǲ2Y���+=ev|?{.��4�7ݍqp�����Ǜs|�e�0���@nt����v!�7��^4P�!�����I��#�>[�������� ��W[�«.����5;�1k_#V��9Qտf �<�i��UvO	�ug�:��(�}s��ꕧ�����y⤔eI���?�M�j���f�ѭP���W[��]����00��w*ż�VXڬR.��U �����\a��$�Q����	��Os;��
va��pʻ̣_{�Ao�mei�.�[�F����hﹴ�����5`�=)��kG:��.�TX!؋i�k��!�e	s]v����X�&����,-�cCC���{�j��C����)Ɯ��,5����?�#����ߊ(���\�n>^����A��ϥ�˄�>V���ꈆ4[%W&o�G�����96_��)�v̋9��L^��Ϙ25���?����g�~H�?����N�y�e�3$n�x��6V����9J>�5��]j:5�,��Q����k' �m�R���Ä1%�Vä1A`H�$���߼W?F���S�=#�E��W���0��h��5s��s@�Uh�ˡ�>�ŞA�L�I��l����z�Yu��H�#Z�"��cC$��a�fav�)F}ݝ�8�*V����ϻ'�g��Bɗ/bpہJk�!: �զ�_����D��]m����̽6ei�����bp�iP����[L\�5���L���%�J7BF,�.ǚ��ԉŌ[%<W/s��աS��ZY�́�{���Z�s.��ɯI�Wv�������t$Z�cĽ>�~�!�m˽K�bӀ��;0L2��F����1�v��sh���۹�P�ҖYc��R�ڰ\������w:�	����n�[���ug�zm�u(�M1`2䐇�����I���F�E�17�����[�]��ϤEDB�q	Ib�A��1��-<��)��KH��x"��N�D�L�yLgO71:%N��-�-�$��2���;�W��9��X";����UO��<�s�x��-n[���M��S��P�F�4�i�+��8z���.�Dc��W4�Z��(H�-_j����:�~�@n͗���:�����[�7��03h���վ�˷����1�Q��q�����,<�ؙ�Щ\ >���ޠ|k0�"��jXVoV�e�a�,X�!�8��.W,�J!�Vo���QK�9c(S��4q�ӫڡ�ܳ������@ˎ03�`�ֽ��T
'Mc��Pы�8پn��h�1��8	�[�\����0:(G���o[�
��g��{_���^T��c�Gf��r{fC��w��(���tT����Vj���i�i�OK��.N��N�(� ��pޓ}K�����8[��LWD*�f~�,Jh�� �N4�k�i+ O}�&���M �s�﹛���T����N����]�oHiUZ]d#;�.��#���U���ԓ7��	ZT�QH}a��b�%�����H�w尦�d�EM_q�g@@�%����o�͌{u��	���v�3�����54KA���U�0�l���TJ�]����M)!��i��p�k��GnS8^��\�:��u-WD�`
�����BCRh?I0�%ui��t
e����֪H4�,.�a[�(�3/U*��Uhy
�%�BzuXJXWU7�_� (p�T�i��J��
j6��j����*�d�b=h(�q�.�!�
msخo%|�ݘSd�a	W>�*Z�e��WG�^��p=gH}��/���'ks�!�eC�R���)��f�I汈o�-�Ci7+�MC�w����ю��b��M~�.�"�oǕ/̘��w1�}v�ވZ˼�~�bi2>��K2ްLh=��F5^��~ʮ�z��%�s5@s"w�N����M����2.�)�	�f�a������[�������,������46/�X�{�X
5��qOz���u�����}��P��f��sA�����y	K���EL�((�Z�#FT�#+����O�٥E؈Z?�����%���X�)4���!vl#����*ɕ���֠�V�ɢT�m�p��L$~h���P�9��[���Rb|Z��w�����tK;v'k�;9�B>z�&�.ZVa�kr�CJ#���{qy\�&�IbK>hw���)���j��QB/��o"�Y7�T��^�����{��\ej�ZYXK��*����pr�N~1!�e�σ������" �K�;�7�ϯ՗��,ԍE�O^ap��s"qyJ�N�z�?�]��&J\�Dj�2P��X�'��!�!QIgR�m��Y{xG.K�n�:Wk���c�� �'��wQ���(�Ux�tt��;���D1/�j�)�
Ad���E\ĭ;K�N�t ��Φ�wڄ@o�����_f�t���sV2V���<������]�� �"x�y�vzd�
[*V݂�x��GH_��*�����؆69l"?"+�����:m�a�OX�RO�����z��;و���]�@"�ϔ�ns��p	��!��h�� �1�#�qP;��V��~/�����#�;�V5�=r��.��1�]D��X���!ϴ��: C<���~���z�ԕKJIw:G���J�gfl�g���$؛Ҧ)�jȱ�#��E�{�9��U�V�&BH�|*����J4e@~O<�%3���k����W�%z�I���o����Oo6B����'�E]�!Ο	
�����R@a�D���7WdO��=Y��{4.[�K�XU����v��e�cs)Ԭ���cͽ�����G墆f �Q9��\�!��v��3����i���.F;Pȓ'��+?+��	B�Z8�>u�#"w�xr�ϭT��U��`P��,Ą�*f��-ZQs,��$��*g�4=��U������h(5E��۸�H��i7��v9>���$���^l�g����Y�2E�V?c�@��R�}�s`��w'����v���g�읎�@x�"\H��ג�y=�h��¹�/2Pİ֕�X;����Ҧ��V�O��>���Ň"z�VHx��\� ������|�>�nm����y�cKjM<��b!1F݂>"t��g}2zVn{����	:��t��ﰙD�Z���N����{����UO����\�,�+z��0�w��{��?����Nj{��_�DsB0A3,�.ﵶ��������N�M�4
'ǟ�Tr!jVN>��i���V���¿�\KsX^��z9���
qd�Z���=@E9�,t�瓩���,�N�5���Ч��cdU��k�!Z����_��ҳgf]Ny�u�����5��7Ҝ����+_n�0���W�L����l<ej��f�F،���8����ޥ�\�XoO��ضzvv�|�3t�w�n�K�.RU��ӷS�8��5�4�(��9�-�N��:�ٔ�@;���c�ə+?2��h��=>�+~D{�ŋ��P��0�ֵ7����*X�h���!�3w�s��ӂ��1q����$'��I��5����9P
	��V��U�IkA�r���g7����}TyGYBm�������N�1[���g��oW�z��/b�8���/�盔���lN��d����foKS��k2
M'��G'�>Ν� [>o_bj��O52,��I7�QBl�i7��	d��x�>g��s��J�;���?�,[��Gz�E�c�M"{6�@��8�ԥ�_[��N�'��^�;b���T��\��G8�N���nه t��O����1�����錰.�Sݜ�?���V�P��qaI��N��_J�ɻ�qo�lS�s=q J�{��������db
8���&��O;��	��䫃%��J����/��w�#3�]�?�~:8��Aܓ^"i촍��'alT��NwG��צ�0��+�1B5S;1clu��k��P	9]��:
���f�I�?��{����6�9nE�_SC�;&�K��Η��~����� ��L�O^F�)������J�J��,N7ZӶ���e���z�9Dw�����1�ͦ_1���D���:|(m�w\�6a%@�Y���w����Ф���ƭ5ȍ����F��.�<����!Gā�g���ݧ�u�xogb�����t�lx�t%���8������ם��g��YY�)��7:�J�Y,�gF3'���j����~meC��U�ף�w8D���{��v�z�-����L��֓}.4,������i=�QDlK����w�ix=�CQ�]��C��/|m���Yb���#�:'̓`b΋��9+�K�u��SΥIL�սp�����y���e
b=`"n������ٰ����]��ݡIlJL����ܘ��G�pD�y�
�+H���=n@C%����,�tt�@~�u�Ĵ�d��1�o�O:)ؠ�d��\�@�!�lFq�r���1<{�o��<vw���H�P<�?K�
(=��ӣk0Pa�:�?��<�7K?@�k�&�iKն�1�\K(LՎ���?:����	*称������Q�F��'�4�G[��Ŵ�KƲ6��0���?{=�rY���'��MQ�ע��`lV�௉-Y�7O�s+儛����wb���� \�ّ���3�'��ৼ�||8�)N���>���a�A�ݶ�ИB=�=�ˎ&��^���Q�A��N^���=HQ�Aٵ��v[�����m`������,j�����J�ҷ���
5��Dy��)ZI������8dn�W�[�,b���v�H]U�X|�wn��~q�A{WDNY6�ҥ��z�	�k��h�@3Lf����
�,12�E��0�}u���6��<��AZ�`6�M��^P���S���R��zS�4�_c8�p��[UAb!6Y��Ȳ��o�Hӳ��J�L�m�0���������P�E��歸�J�Ӂ�Y�3_�U�S06̢=�N�2&ܶ��2
:� ��;5ut��������s|����~��X����:��v�s��}S��ޙ�t��	��#�#����S)��]@+n�sVB�h����;�8j�?Cl���f�<&L��[���6]�)¡���"l��1�殂[��\�vz+�n�6�u�@��Y��U�H#���U�)��([�����,���r+���>�w�� V�`/搟�`OSP��Uc��������*G!$s���<s/���L�ӳ2c �͇��w�9��Δ�df{4a���B�l�O6�ӛ:;��KP�#�C�׈2�n<.7�خQ�)��Ko	��$�1���CD�w�p��:�C��� nN](V���p/�R����n���d�cDC�[+��X:��l��U�4MW����|��ɯ6��bT;����n,��i��a~Ե�\�b���#�f��:��?E�NΧع2��l\�����작��e�_��|�rq*�3$�j��!�&}�o���%���|���B�ϣk� �r����(�����?T7�k��Ҳx)�p��VSP��H[�tzU� �v՗J���?����]ͫxl��P�T�6����hGe��EՍ|:���(��?��Pv�T��jy���d�^����/й�j�;��l6񨗼���vM�ǁ�V�~䔹,�,v��߈$�Qx"�]MP�<A���w��s�+��$m�t>2N�z���L�3Yv�(M�?�苅NR��]^���%ſx@v&�����\�gW�q1��P�'<���}ٖ��Tj,@cy���E�܃ɻ7�`�+_U�����ؙ��r�NU��F�}>L��F����S�!�[�̰��*!Q����3=���X&z��v|��́��E��4àT
V�b��������V-%�dI�B�O����<,@��~8 �2>$Sݺ1�e��"md�+y��Jr�$�Fْ\C/�@��zQ������>�#�.�0'8�.5��:%T�J
�����(����!������٪u0I���!�!+j����2�N>Q5_��-� S2����4ƿ�*:Hbv
������K�cPS���&�N�3Yξp���xN�ń�udf����f[�/���;�&3��L�e�YLԈ8�sz=�ĭ�������;�����\oq�B�u����5�Ľ|�J�6�'�G����7�q��|��6�֏X^1�&����"����*~��vた@�h$3���-����4t ��'�t����wަC|2,�� y��P��!����$�%�][b�U1-���r6����y!�=�.>�F�M~�ţ��Kr��v�<�Ի���P�&>絹��R>Y@��Ů)3�*+R^�!�S��15%�����m�p�g��B��Xek���#��Ih(@qL�	�}YL�F86��2�'io;,s'�*���Mx�-���X���|��[��(�z������쏄����y�iYq5�C�G!́5�{]�"��/�h%����-~�p���r�#�=��Mb^H�XT����bS]՚̈����F:PG��N4cE�O��139l��0��[� 	��(h1;�LS5�q�IT�©&�m��R�=������S[˘�i�i�S�q�|���$���_�k�Nv�!�"�7�Şcd{"4)ةXI��M&����(�B��|=�C�9.��,�%���G��VE�P��L�[���^_6X<ߣ�c�A
t��	�P���(�rwHtVx)�z�`9�����ޙ�5���h��\-��T]�=mW����9c69�֓J�5�	c����$��ۆ}��K����}��m�� y'�R#��`���N.�;����C3'+E���c�_v���q���O!�}j�G�������޺�WtC�t5٘fE��c��$]f�� O"����ӝ�n^n3.�~���2��;hϢ�=��L8X"Y�Չ���/@Z�,n����cI
E,b��d�ɣ}�;�ȟ�?aa�}Ui�G�p���m�(���yW	�LȘ��� �2�?հ-��&��ǂn��G"�"�<II��F���[�I�#��.���ֿ�k:��u͔��ɵ=ڒ�8B�f>���;�93�q�s�O������P����պ�����/��.g+Q��J��ه�;{�c���K\�,�E=��+K�"~Z���J~��� [���j�2P���"ֻ��� �̋�B��Y��
�R�B����G��1|�!R(P�&۴M�f���=��5q�SCL���A1���3~K��#��3fJK�Zwm�CU���os�C��YUx$�/b�PhƍZ����������f>�x�J���!��0���^�_Ǥ��*�A!�%Lw�m_~��%�!w��e-��; ���5?`��s\���& �z$Ȼu��K�+-"�;���;��$��o��׳9u��͹[[��W�<�&�nO�)�� �&�1j=�y�!�g��*�q0�6%��^Q?6ֹfl����v��wT�0�e�7P��]F=#���+]�X ���Z�n�F�C#k���2�ъAa�JQ��5,Le�fT,������]=!�5�Ԏr��Phb�~m���ļ|�u��Y�mHk2���?�CXBd����dir�L�93��AQ�.����o�c�UD��2y�$�{e�Գ{�HVp�����Tn���{�İ?lFs�d��QϯK��g��ٽ�����{Q�����)�f�s�s�,LJ�U[�%���bQ���'D2 h�#�}���@>�/�IpMۂΦ�;Ă��S�R�P4�I�J�\��4�/g+�o��!j5�c�r��M�t�Ǵ猔���ʇև!Y3�<�����9��\_]X>*޼�(x�_�V!�%]j[p쭇T7��.6>��"��P��`�Z�>���
P]��D{�l o!M?1�嚰��)�d���B5 Bb.����
����
}����<0B����>E
K��@�C׹�MgضS�r�a%��뫈^��C&匠R\ܹ��b2���ԛ^�O`�����i�e�;P���u��g/�H"?2\�ö�b������)��0y�p���k�)5�ވۖh]�'o����Ϸ��m�^\��j!+�,Bu$�s�Or+pf�6�?U����C�i���� �7��q��u�No��\�[-p&O��/��ܴV� ��� ���o�V>�X����R �k���Е�e�N�Xd֘c�L�.��	X��^��)��*�������Z{��]�.�`�6̾�?%4C��ؠ��A!���Һ56:�"q ��Oٞ�� �w����"��Ez�{����b���@���B�RT|de`����� g�� 9����k����;�h+l��A�Rأ��g������7�=��&�Y���br>�[@��Ÿ���h��y��gZ�y�$Z��2�^���^�|�wl�X�3�p�M.����4OJ��BM�����[N?�>�<��VQ%'4��YڹT�TFo�!%�	Na����%k���-�ީl�� f��X}+گtB^��X>���L�{�Ǡ�=�7���T�N���pC�Oa݄#�ƳJ����24w)[���5o˗)��e=�)Z1'���h��C�/�m(�6�K�>��4�]7��`k{�%�c�L��H�hk@��Y��`n�y�G>�k�;�Q#d;��a�ݩ\��,<�٘UIzs��m�	���_�߇>�%��uws���]�ƕ�[�A�9T��h-����B�̬\9����{ʿ> \G(� ]t!�[�xti��Z���������CZa[:&���vi��Q���3��	X϶w"�O�z�����֜7��'��x(�^J=0y��%��&�J~��k��H.�t�<��S�T��$��P�b>C����ɎH����6�"��n�%pqqVU��t�{��P�O�Bb�h�����MI_�W���p�`�Et���ñ���a�o���I
g�H��v�.%/��5�]k�҆l���\�Ů��]׽�ŕ�~�C�y<�y�6VH�PhN8s��^844c�%R(py#zA�D��$��h6˙yX�."���5���ҷ�S���1a��2V�=9'7�4�}j�K�	T��n&�n���޷�m��.�j����ۥy6�g���69�W���{�f�����ѡ����X��{4�3��;���:�C�`��`\�0��8�����$Dz��'�P��BW�/���b��m�\�$��Z�ֿ�m�C���*Z�ch�G-lo56�{��7�0��u��.*R�D}�\�}(���B�ꮆ7%�Q��7��3ᵨv@"�t� ��E���>Ϸc�Ohe��{�W��*��gM�h"%�2����o�:�
`�1��3�-�'[�R!j��!O��7�̒y����4�
Q��i�,֦*�2��L�e@�+l��@���V���`
��%4�}�; T�{N!�4{\԰�d��<��u��θ��ݪ�E�v�P���{*���n��X^�"z�-0r�-�����	Z��<ؽ��!jc�y>�j@�'�|�* ���4�}	�#���m�	�NX'�9�H7�t'Ӷg[���� �gg>n�?������i/i��RSb%;��|cX}��`s����g3�����ܟ��Z���#^�49���Fl
E��{����g��#ma�=�rԥ���=޺ηH��~�inG�'���P�Z�W.,�[錯�֑z��]ur9v��nk�b����~��M=7H���ցV�a�ѿP��t6��j���������3��b���.�ζ14�fn	q�iS��ó��x���,j\/G�8��!g��)V)���⺚��Lq+CR�+Hw�����BzQ�"�T��(#VQ�j�T?eK@g?O�%[+�p��B�pZ"�:$�r�N ���m�(����8����z�Y����hA��=���MX"{��2�ź�w8
������� B��� �di���c�	��5%ZF�ƥ���2�͙�]g��I�P �����������J�Ɠ=���<F�%
lzK�9��]�=UԂR��]!@V]+k�G��:��:��A��ɕ;u��J��Q��$�]�/��1��'G�B��/h5�Q��G-O��G��(_������Ka���%��B�O��_7�3��y���}nu����sm�76fI�x)��U�kX03�t��p�؃=	�bvk��9���5sTJ���� d+τF:Μ`s��c(1��Mm��D9�t���u�?jOqy�M�|����d��%m�h2q�\��o���6���o����ǩ��]�"�<�����(�O�H'ox]�����#+<��mb@[{ދVχ��'R� �\�c���̿�)[q��vi�`�ӕ���*�z;�Y���nw��}�h|Q%0�|�Th��jk-��}�[����Pm)|"�Fc�A��w���v�UED��-;�	���C��u����=@I��&SW������#xA#~ЀI��Y+���M�{٣�7V2l�
�Z˨Vt�-�������#0�fH��T������D*͗#H�A����O�W��4`KSF�����`bno��뀢<t�-D�-���Y�P�����}_g5>0�`Tm���8�����I_��O�<��h��}+��-x-��,ɛ�$r ����qs�~?�/�Ec����IM~F*�����x�� ���
r�z�U��N�\������S�@x��+�=��>������#~�xz�kx��҇�G�kB��4�Zd1�?��������gǵ��2�<�{�qz��s��$NwH���p��n�t8�@`��ؘ���O��FR�)�2�.�]Fb�.-�2�>
�o�*U*�%2~��N�'ma*�p|��F��q����ؚ��<�_A�B�p����ʧ�mf�F��5���"�\b���YH>�N�!/�ge�N�R��BT����g;�\�MF��0f6&��s)��v�)2�q�nf9K�4��T3#&��q��lcL����i��UK�љIM���Om�e�"8�?{ 8�!v�Xi[�eh��xq᫶YQ�n$�Zq��OJ��U��\�ȇ32Mxl�:/�� �A䡗(�֛We�p��:��Ha���q|i�� �ɰ[QP�Ŋ��р�����%@U�Cr7�5��̽֊�<�,R�(��T^�5%Ġ&�H���'(�B�6��{�i�F��Nb|�Iî�Aˊ����s�j�@�R����x�
�T��+����-m�]o]ʮ�5ޤ�����9<�8�jأ�L.	:H��$����e؎v�ۗ��ڄ���ʷ�l�aN�g��M�Ψ8Ѭ/0E���XΌ�a�4#bc�%���s�r�65��Tx/��m��Q�N�pq�D���������,B���=p�.ӂL	�<8ue&�X������H9J&=��ͱ���Ӧ�Ў�Y�@S�,w��\-Nu���.�h`��h��$�R�6p�n),��U��"̺dvT��]@��y+��T�k?��6Y��p�x�}��\Ly��"4��Q{�O(r������PL��e�;Ϥ���=�߲���7#�t��EI�[N�dľ��Q�Uz���w�u���*�iT�T���w�;�.�����[��!��-��T�k����	�3��e���_�+o*�.P-��R��<��~V`6������$W�$���M?H$�躴��F�e��#{<��!��%p*:�A��Z!��h
�vq$�ĥ��I]mE�3vLV�&/|������r&�d\�%6eA�M�zP�`���_s�U�풕�A�A��:6��)�����h�!�{�	:�������'�����_W"4�x؞�-F#����4�m��H��F�OG �}�WP$��_ԂDQِ�h�5s_@(_&��٭x�S��vrjL�����9Ə�MUb>=��q0k�5&�
\�e�E�ސ�:���!Q~���WD��1�b;ߖ�R�`�C{C?Gj�������)���Q�����s��Z�J���6:4�YAx�ӡ�ۯ�aΗSr��'T��������~�#�M�^wא끷�%��Xcc��X��RSl�-1ߡ; �BJZyYR���Cx�ͽ�F�\5~s�8h����a�'���ʜ���V��9=��!_��u���qҊ�m�c��M��̪C�1 5�C0�B=�~4����l�F7M�,fw�"�cn5��HqUх�$��6��r�^z(Z�?mx����L�\FiD��[pV�D��9�&�����	ܐ�����LXj��Ŧy;��9����9�G���lK���Z�v�_�<����&2i*ߍ�|��"�������HG��۞/�@_xl�#��[owRx���?�m��^���4\�h�p�Rf��t��1��?k��=I��ِ���G�j�w�Y-7��Y�\����I$1������;�M�S+.�YeZp�I%<��f��2N�����$y:�p�8�V��Ȁ�q�y�r���s�Y�!^��8���F(K�0f= �����7%��p�G�陈�e��wb�v;c	���8�;^��02�-2���`HO��5�F��L$����o9%��R��r�w'�ԴPu,��H����Ϣ�z���p���/��θv��}�;�s�"a���)���)�J��cm���6�<�p�J���s�B�ԑ�D�X$ݬ��t�L3>i+�ۂ$a�xںK�bf;Tv��OM9�hQ�D�U���P��_�6l9�l���4�5��z7<�\N�ҎS���1."9��k��K�q���D�:g>��k���Q
 �N
�<~��%���*mwq!~R�I��]��.��<kh��7K��V���b2��A��oDN�v��L�PA���ɉ��.9'�5�u��,�BpԚ�A;����
�+�������l�2V�%;��8�|��2��vx�K;qԾ�&�[D��r�ͬ/nU�B �E�RX�`���Jv�s��M��̰ ��9�B��U�ފkYܢK�RA��f)���v�fHw�����VO��|�:�쀺���s�����z�'����HL4�3׺Dk��g�+���j�̓�;`�T1*,*��'�����ͅ�.K��0"��(� �r���^u�xΜ}���|�)$i���)��>�$^��o{~���6���?�f�m� ���X�)�$�5-;ܬ�W.�|��$�g�]�Gi���6���l ��8IM�w�"X��6i���C5�6P죘� ������Oc���˳Qa �q���\���j괔���PW�d�'|�SX�'���JA��-?���ў|ft���Z��=��mtf��)d�A������"dAe��%�z��g�z����D��2��Q�[>�!g�-��&���O�otb���m�(E�%r%��Vt��M;tǹH{�B���	Om濁HY4U4���s'>���<"�ДY���S� +v��sR[4(���-�v��	�Nɿ!K;z&ld��#�i�*�]��-���;�%������4�����F�[�V��;��&ׄ'!f#�����)u����1��K���s����&E@g���/&kL�ϞC/EW��@^T�N��q_��� �LG01��i���s�uG�Pd֞7~%�婝��9��Yc���Ib�k�~q9i�6��
~EޢS���2&��=1��Ю�
�P��6��ak����:���H2���>T+�b��x�r���F5I���+�<���/�.�;�O��ԙQ9�.T?i`|$�ܢÁpb�W8niߜ�'�	
�;3�%f�c}j ����&BvMr�޾��MǦ�)�d��B�ˏ�������4���-�.�s��Ä<�4�c1$�"f���G����Lf|��2yt�t�{t���CYP#���R�^��lGx���Ƹ-q�M}B�ĵ�~C �2�YF1e\=�����o�~�$�4d㽺�:�E���b�\�xD�J��A��;�P�
1�F,��WYܿKPf��y���[���s��p�W�3���fc�H{ �P	�
�B]Q:̱����:_\��O
8���ն��0�U�{p������L�w�O��������t��3�pV�e�=���X8hq�'�]E� ��	��n�	͂+(�$�>���}]њ۪x�����c��Bb�>�F��[��dW��ת�K�4��M������ͻ���Gk�c"_��5zS���ї��v�7��^�h��[8e?���[�G���s#���,m��&�e#��m޵��;Vx�������޿2}�&�l��P_¦^�źXe�@]��K�����X]�5E�S/o�5,���h!�~&�;A�{/cv��iLȅ��;�%�k�5��������ahz�?!�hk��t��.��}��{i�k_]#��q����զ㽺r^9E 0fY{��h��W�;5yTF�h�����ai�8
ӵ���sS�U�򫜁�K
��`��<|�����ޚ�yѶg%V��ڰ��}�Mv�L��ep��fr��ڀ=+�� ����4jP������ޞ��[���v��ה�b�h�U)�p_��;FA|�B9��_��k���Y�
%�Y���-�M�AP��b���3�k@�ɥ��I��a�AR,��:���ä��� i��b{`=�֊��@�uq�3��}�G'���z����婥�4>�+�����	\}���Yd��4�� �3�{T��n���l�u���iu�#J�9�$B0ܪD}Yeˋ����j��c��"��Bx�xg�<��m��[+�.���&���ҡ7�M��3;}���k��F�`�xP��r���l��v����s/7��ZKTNV�B�$ƛ�>Oy�׼w)?�RN/>��;A�LZ��[n�tax0�3*��u̏Y�e��%��T�G���ycTx W����œ �����~�7^�I��I����]��6��3�\>�I�l�/�:�F'h�b�O���ΤZ+*o�s9J��uj]�;;����
�u�q��%B����z�A��M4O}ʱ�6�EE�3B�t�������n��B[����A���`>J�������I`.GR�Q���X2��q�7�r�X�ak�N��%��T[��$|M&�� n�I�~n�p,�p�q����P"�M��pyc���H���e���d���*�4/W�_Tb=A��#����)(KT�t�X o�w v��C����$�K� ���u�w��떞�&
���i�r��+�{F2<Oe}�����6��
Z��g/��R�#!�\�,:6!B�t]�)���?��F)Uׯ������z��&���-8S`��u:��G��I�b�5�#Ρ�q��}��*L2h{�5�3tVs%�d�%@y2���l����9�aeĔ����'���N�Ȱ.80<gv��O22��ꔍ�d?F�叹��V�+�4_v?C>�k$��w�pr�:(���+�na�����/��~l>Î]�������q8;�q�o�6�8���5�HV1�b(�)΄M�����n��?S��z�la�L�X�ah$n뇸�ghi.�+�y�"��D�S��;��1ʄ$���2�ѷ�`��d,n��a� ����(�$��r���U �tZ(�����뜆�j��^�l�b��f��cВ4Њ�U~v��S��c��C$`?xՙ��ݑ��h�+�ъ%��Z�N]��'Ň����X�泧���a����?�#��U�l�xl�"����QBCx.�/��SU�JP+B�OO ٝ�A�س�U��.;�E�j�+k�.}����N�����?P&�W�6��<�=�R����ͅs0�.qjh��I�=����B8K�M�����Mp�-�0��ҋ@~C8f�5L6.�6�H#��y��,}���Q���u:VI������'��� M�Q]�6�)W� A%GK�j�}&�&���t緀^\锅���J]N�|:e�J�w\�\�B�1�,b���䌨l��XT���>��g��NE1�j׸P4����X�c�]2��+�X'�B���&�L;^�_j_�߂L$�������}�g���[��i���ݪ��E�m��F����-ѡI����K1^Ȑ��6J$���Tg����j@��tA⯗(�_u0��_��Vb��^� ��iL��SD��r{���\ﶁ���l���f�ޥ��1�d�#���iw��ȂF\�'���k��҅�g��|��e�Ӫ��`���+�G5�j����3�I��-�-�)&�y�f�a�X�?)����_���nHiD�b7FMg�&�V���j�¸<ގ"�fP���!^����{'�Ϋqs!�z!�(�Ƙ������'��`s)mR�Q�-��%N#��� ��^ĵ�ؠU�Rы�U3w
���$/��at�2�G���������[|�q�n���ޣ�CN9/�e�P�E�U���J陂�:�0�y�k��=9����N���|{Ժ ���G��{R�(]�S���?D�8���0�t���o�ɖ�����J(Y���B����.מ@s����ȕ�?0#E,�̰�l:ib�Ca�!�Rٞ�)�8i0D߻ښ%���� t���x�e~�1���i���_q/dQ ��֍���+���O���BӨ{��W��"內ER�I�(ѫ�qs���ˀ! NV��C9^Q�	yb�a�: �G�g��Þ�1���ң�B������G��C��ǟ�s�|�����SL�y�f�.��NhЭZ؝#^�}�H��~��U)���L�us�(���8�:&���ә��xKx����1j���<ҩ�|p����<X�)�1�Q�hJ|"�˼�+<G��oee���?,e'S_�-��0v����^�7taΎ����tF��!`,o�!k�?��T���nb�1�\�N����x�����&,�K%��N��q�{
���Nj ~Іd(�&���?	% Z�!ʁ1V���vh�־+[���e��B�1�<T��e����;m�QEO[��ӊ�[nl��RW�`��cL�qrz��a��i��L��Y�������I��	7�����f>J󧚵�_f��o���	
`<Q��c%�!�-�p=���͙�nN�~^��[�B^(�r�b��E�v�4g��fO��{���fW�8%:'tP�t�

�A�~�MG��o[?�I�T`5F���ydh�Ö.ÏB�e[k�݈%�k0_x��}���N;�ԁ���Ty�p�2D �~9&c �ۍnfG̘�i"��/�F��,�G�R�U�P,�!W\9�`�\� XC|��<��ۆ�[��|W���r�}̰9�̓K�f䠘`*P�>�:Q���1�s��>l;�t���nQ�*<_9������v��{��C?����@j�$5$1��+�tQq���4�	�3�a��)ICu����(���TpmIq�O�����-6B�,=�U�h��>�բ��E*��ڵ���2���ϵ?��V<�M
���w�T{Z��/w��?kг��4X� ����Le��vJ�	�vZe\w���?�.D�D��р���6��Q]Ħ�TI���)_���ƕe��7ʰ-C'�_޶�f�˯ʇv�K���*�����A0I��?k��[l��2�X�x�A�|���-f�q�*��q��ޖԋ  l�ʉ�[� ��t�mZ�}�]6ʝ�W�j�CH�q�"�f!:�!���}Um���<�A�]a���QV/�]U�rj��xᓘ�'2s!e�4�Xw�iűqVs�~�~8��'Dmn_ɫ����c�Ul�Fg�F#
��M�aO�%߭1Ĥ�s���|r*:�'��o����-��%�b09���Evz�M���*�}���]�Y@\��1s��P�ۅ)��T�A	��o�O����ef<�n���;%T>%/�	��DH��ө=K�ߏ��tr���,=b:�`<	�]x�����B���X�_T���p����������A�k	�^<�i�I)�{S;�n�kÍ���`��7߷y�v���7>l�ne���'��0�?|�}��eDBR�z?4�+�	�����Maa�k�J�fW��n�'��#5V�89C;�+�1Lh�kx��ʞ��]������4��'�*2��
�p�:���ݢ���z�YPHKś�m�9@.�T%��p�߄�N�y��xQKe�<�}� B�]��&�j��;x.�7å�}X3*�G��Wh�Z�f&�J�\Z�$N'���5�5:����ʽ]�a4������O&&[�z���|�z���u��$k�d%i`�bp������dUxK70�~!�h���y�5��u�V�����-������nS+<@M��%����faZ��X�ʞ�EO4su[O��W�]�'�AxŌ��l��� �\�s�ٗ$��,����h)\��ދA2�gV��"���>���qxc��"8��6+*��;w�w�U� ��L��z��y1�n�E�8mވ�L��~䨆:��DKR�������?��W~�ԌE�~��l������%!�;ӷ��G�/k�yb��_���H2 I��E�j}�w��[�����C�wi�� ��!o�#�W7�¾�嗾0�:�	?͘v�S�N|�<���a�����wVvsH��k�b4Zq��ږ}%Q<�a�g���7E ���i�K��U���vo!,o?iя'����������V?e��ia���}� ��T%D�fCY3�:�֯棈�,��/]�4)i* ������u�ʊ'�a���"�x���m� V@�e4"��ixn?���J�)W�Э"��/�8�����e��+�6������F���ǰc�;��4F�C0����o���B`�%3:��Ui���H��*yN���&R,`�`�g/��^�@&��߽Y<~��K'����՗����\�c@�ي�.(T.fkՅ3Ր���6=ɰ�A����]8^�:9E�zH��Fy%�h������\�8���a�sK?��#ޣ�����t�b�	��7��;�Mj�6�`�%ҤD�I�I����Y�I��rf<���Y9�I���k��"���z��*5��T�	�N��6�?�֕'~f�o&���	al27�A��������+���
!{ �ʇ�g���{Љ�R�Oqo-�M��7�=��	� f	ş�X��Ӏ!�㕗E:UM��_4߄c����O��&_�o>7[�"�$Gx�غû�]�� e����q����D�^��V)�Q���=����k�&�7�c#����$�p�oD��<.�'�sq%��PW�'a���{�����D�'L�qj�˔{Jˤ�S<>�*m����q���!ǟ���F� >/�q�h��Ѳ��$�S�Y�~��Jf�ЍN�,l1���O����q�"��7&��c���>M�ܿV���7�mr�!t����lM:Y*!h��E.Q���I�YsE���V��9��9@ޒտФ탃P��G���u�)u��y,{�Rǧ���M9���_Hx=ҿ?wv�g�E���o�S�]O�����jPb��Azѐb��L�n(Rz�U笹%?�OK�Ӵ�9�]iʎ�b���Ϥ��k�;䜟s��L�+r��g�Dct=�q�K���*�(�v�
S�$�|iۂM�$ll�q8�y������1E*q�Ő��w1������wZ?!Āt�>�Ʊ�>�X���(���g@9�����L�(�B������h��*w�# +&�ޤ60��y�Ϭ��7 p��I�Q9]گ�J��#S��%�_��Wj��LiCxW�b���qr�b�㡆�v�!��������tRb5�s���[�,.O��V+��]�E�"4(5Nȑs�\�i���ϼ�J_ܴ޴I�0!M�j" ��Ucg�M�8��"���F	nN��3ԍN�z �񑏅��� ���UDs(��߅q5�a(@�)�&nUc�+�j������u�%ᝇ�NV`ob��.�u6M��������]7HƊB�
��1���ɀ�P��k���9Y��5�h'\-�ELʠ�L�� i�.�^?yy|�B*_��.w�7]�)�6(pYx�h_��Xme/�d�����=>�t�� ����>�Xp�s���IN �UF/B����m<�ҭ��e��vO�P ]h
�����P��b�U��.�W���V8��D���Ү�q�*�58"}\�F��_D�T��q�q��6>�%r�0��N),,�U����%�� ���u�(o�ġ��8]p+� ��K�7$5�j��(�-���*3A��K�ߩ�t�b3�ة���ԷQ�����k�F�\�v��:���W���Q��_��.x�<�,��b���%�l��N��N(�Q����m��2��u(	
2�cg9 �nH�>l�g�2�A��H�&��D��¢'M �Ѡ�g�����=��@��d�Qbh��y��-�)k��QC}46´&��P�I�Pv�	m@�T��]P��鿢�s^��9=����ۆY���;);��_�I�8o+�KZ���?+�X�ZFN"��u�T�P$I�m`�)�Rx��.�b��\Waq�B��1ۄ[&��~|���I ����y{���
���Kf" ��U8���D	�<��n!�T����%L.^
xC�W�r����ǌ�!{���w6)���j[q��1i���L
��,?��!.Hl�l|�y��g�v�8���gG�Ek�C�Y�ڏO���^�|��`h�7�V� i2���/;V8�$�v�)Z/�>�mC�����)����D�e��� pnr"C�'��;��7k���~!x�)�]��͢�Z���͎�+�`�T~���c>^{.W�R�)��SXb� �H�hΝ���wg3xRQi�>mn��&�h,F��懱�ي�����J��U��N.�*�����t�p�Nҙ��x�
C["}	^��r@�h���*J�`�� ^����e�p�s�@!�6�rƫ0% �=k����Q��q*���P��%�4X��_�<<%�1�M��2X�)�I^X���f��rNh?�냁��3�e?�!��h{>�������UR�Nٱ>c` ��a+���	��?�ٚ�f�	��S+�K1�w6�L�:\��{�O��6�7.�@�/�RH����Jp��w�)Η7(�|C
ӿG��P�$g��?�{�(�ߜ�sg;I���6U�x�ة�o�UWD�?\�ͅ�v��Nk�`��P`�3��c���X���}h�N��,��Ƭ�Q�1�3Q^�������薟�kTq�T%�����4Z��9q
��-�&��pk�k��nU�B��A@^qo�E��%�`��*7���D�C�yc�Wn]�Nm[��^s��b\`��I�u�,�z�Ԯ'V�S�b8$n�8LP�� P�_R��s��h�'�k����=Q�V�+��Ҥ��;q���G����ivLG���4�<� .��4��m'��L@sŖ����4�X)i�һ*3$��(�&DQ?���ESn{m�٘�������J�_L?�XuL�G;\�U7K`���.���3�9�fU�Me����ؓ%����*��~������o���K����u�5ļ�2�=�.����ʉfI���R7	չ�pGт��D��ϐ�V��}q���w�8���GR[�Fi�g/�~9�NF�@j�z��5+������%�~N�b=˹�����z�M�t�z��ς���9c_� �^�9��IÙv���i����Wʇ/�$�d��:\f�jn��6�����9�=�۝�@<�`�,w�W��t[βvzwy�~��=Ϯ�s�v!�����zʺUn\��7�ڕ������e�(?�4�m��~�'�s�� ����O�xU���L� (t�Ce�DU���V
-��rGM����g��L>��<��$���0�wB�3�_<?�[
�Y���6C��ɝ:��`h��p����4�\;� �����~�DM�N&��N����>¿�&U��n��� �w�sGV����"���' 5����r�FD5OM���i�N`�ł|�%���%�H���W�g�ֿ%2�P_� R�|�"q9B0(��KTH!��pw�x��LC��'�k@E��@�gQ{�m��B��~հ�79>@_v��G^�œ��oL�A�Lj�^�?��dM�r��QP]P��# μ!�0��H��)bl��_Ͻ�Ś���z3�޻Z)R�
�{D��;{��0�)�s�)�$X�j�pܯ0���Sd�E��ditj��r���&�����pqW5�b�wژ��N۹d�^��{cȥ}s��'� n�P+���m#��� �:����[I �H�?-ie�T2�YKtI������e1����Y���e$��-%)Q�G�%�}���>�*�p����ٝ�h����\h��F-E�\'tE?�%d�ن�T>Er�h�?�R�ꊈ���o�n
x1���f&��k�si6����r��^���)�NV��o5���;񨅓������=����5���'+S���OەF��*�VM�?rC�ϧm'���A�+�1�8nsg�e��Y9c�P���jIL�5�����P>$�׆��lMV���U�h�yL\io��f��;)k��6�L^��Cס���n�z؉Z�����xD:&U3�g������~nz�~b�ۈ�if_5}~|!2}�1�5~��k4�M�q�N��s�3�s#�� c}~�^���i��@�tډ~��e�\#wʊ?d�&O��ǱYC���\'�m�8�d��� ���� ]�����Y Kb�W���v�\c=�{��䤈�o�_�.K�����FG �9d�np��JO��Y"\�������� /�Lox��7;�`zLl`�dh��p�������uѠ~\OoɎ�K���~��S��#Vx�/�v��&J'x�jF�C��\\
�I���o�T���9�#�u3M�R?�L"�Ds��MU�r���&�F������+<b�@$���
��N.�_��Q������p(��Z��Xë4�x���S�ґ*�B����T�bDm�,�2+F.lhM��K������ȵ�=6���9/2��u�^��{�����~띤�I���O/U�烪PhVzB�)�0��i�*Ts�r*����i#�8���1����,jr?v�����	A3��,ӕB�gQ��"�6��o0�D�\�����/�p�pʳI���2!T��X�H��+��-�B�p���]w�#>�`�܋� �M���FqF!�!�������xr������g��xdX��j�U_�|�����#$�q���M��o��s���ۼl���n��@��nVfeT`����I��5�Re�N�9eĲ4�.��@_�d8Y ͏������4c��6�Ȋ����嗽R,�Ya�禕`k���^��+���L��KJ$��SH�uG��
h����e�0�/_4\�఻�ge���-���V���2PvU��q�9�x��R�*)�A�:A��5<mTCK�v���bQU2:�c����ܺ֤�`�4��e##C\m�
Kn>4񇙽�������Y��`��d�'5-#��mL�ۛ�!�V��Y`
s8���"�������
UT����5�rNjuAj�d+��+1e<2m�Z�1Qv�����Y�ɽ�/T�b�X8������ J��$�;��":Q�	ڛ��a6I����͸�}��
}y ȸ�*҂
a@4!�f�Li(2�N�x'��q�/2�e�`�t]Ě�B�	טj��8��{���lq�UbҨX�(��eFE��Ѯg�C{K�P�fW3�[�v�`��iZ�TFH��!CW�����ڙ���4����~��A2�C~1/
�q�_d4�e)��[H)Sh�}@��!��Qѣ9���h�A�m���3i�]�x[w|�V5�sT�L�u޷7ﾉ��Bº��@�d9^VڦF��9���1�4^
��i��-A+-Y��e�{ߞ�����րB�z�s�8M)uR��(�X�)�����ړ1i��Y���vP�U.��K�Q[,p��Dc�0����o\R��`K&Y!�+��r�O���]���"��2����܁��x��L�~�V{���r�V-"��m���9#(ES�e}������cÔsQ%��;F����,͍%Us�9����:���X��T6�J��D�k�����|8�ܘ7Hq|���O�8��=Η�?��p�z�}�޲��̺��A��ݓ�6hhA�ӌ��gi�cE2�����%r�eW��V�{�l:̪d9��=�}��e��9��v�8�`�L} �A�[����Q��RU�{�
�'����^�5�hԬ����O*�K����YI"�I�����ޓ(ʗ����w�v�5��KW<����'��R�f�Nܯ0Wk&�W���ҕ��Wԉ؟��s �0�1bt$�<�u�m*��/�X�G7G��9�(��h��4�������z�FwN��u�_{OT���),�Cڃ]�[Y;H�ya%��Ƌ��[l�S�[���/�Yu�T%##��c��z`��?i�v,���^'�H��=1�>% <?��O,uh��l���w���֛ʰ����X�����N~YXټ Lfà;{�!"�:��nW}LI�g��Y��`��1� ��Lѥ��ٌ*)q��+u{���S��Ԥ������p`E����
d�<����J7�����M�y��X	1)�4�:Ut+��M�N;�z:S�9+x[jb�������h<�Jt�����	�X�poC�h٧�^�+�g��,tY�����nD$�gF��!���ytW˳WNT�N�&@��pC�>�c�O��	,�.�!��޲.�p����L���j��p����U��W�~�k�|�=�@�A-t��O�$���A��꺒<��z��tB O��[��d^��*�m�13.:���>��x�n=�2��G�8��j~�˝$`��2�˞&���R~0ߜ@2@���������k��������4@%&�*�T��n��WIT[�2��POeV(d��=n�b�r��\١��	�Ӂ~Bg���'sl+�<�V�������E�y�{'z�VJ��� �B�N�3$[����d���<�����T�&Uf�r}�]*�X� 6C��UXv�Q���ۺ̶��
 �r�S<h���_��*��}�F�'�W�Cu��4����3?g!T����_!R����C]�ew/�|��bU'.�1�S!�iWҠ%%i%C�!~���,~�C��-�X�zG�겳�&+����K>Cn�,�0^�ó/�+G��,MH{Gf{HnQ�Lb�n~6�J���b'*8�2���&'�,o��g�BhX>��FD$ȸ?��]�x.�rSz���"��a`'���{���=����+�Q��k@�y�otY�6�yا>�e�*�q�Y��w}��R8�+Ƥ<��2�zx�'�|���!���+I�~Ż֥� �9��B8=���a_;�`�̻;g�����R��O;���{��q#����E��O���^(�������,��^6A1�e�mזd&g�u]o�����~	����1˩�ŕe�
:t��êQߕ�6�L&�p��p��ui��xT����-�� �Y��{����p����q$����8��5�q���]�RF[�*	�����<ZpY��H��%m�*�DT���
�N�{+�$8�EK@�!�2Gv��:�>�c+�՜�.D���G�M��.2�A��m*V^	���@�ϱ�9���F���G��#��]����N��˟c����n䨊Rw��N	�燳3Y7yK�&�}� �_AB&I>F�l�'�0�o���D��%��ur+��2�������mr���5W*�����F��.�����#��}��]L	��TrL��l�Y��Q �pmzU��N]{�w�hg�]T7x��<�#0�Ƭ���D�a�M��Kq���i!/duHa���U�]D����~�U�VJ�F�:����m(%�>EO����l�D�5J&��)�>��4#t1U�Ǆ�TX����gRbZ�~mK��U|�~3d�l�u�������������!�FB��7�;H�{c�i���
Q1�u�b*�J.T���D�ȗ�u�LT���:�a} �o_��iZT^��B�����vUk���n��'�8�X~;D��$��k!�v� ���f/J�n��~|S�b���ܫ���:���/��<B��O�f���������>���zHmB	��x���n�ư1�Ƀ�ܞ��������::�Hj�^%�Ʌ0,=�K�"����
�����
�&L�DUau[�������5}�ƫ� $���^䳨�1�eТ�̣nX"G����DIp*�y-�s���3��N��SW��5@b���,�:O5�y1����]�!(C�����c�r(�#���-m	�
8�E{���9V���V�XK����S�L�ʻdIF����^���;��m�	ÅRk��m��F�o��zhnF���9#�6X�N�`�//��O��:~/�M���qE�d����*�����l��/̌t�$C���G ���(���L�4;삉tO���-��Y�(i;YN���P���0G��E��(F�PXb�,���y� ַ���&�)����8Dm������`�rJ�j��s?��~*��q�Xf����h���:�3���i��/l�S�� �i$r��
[�*��J�r��[b9z���"�������蓂���.�?��e�ʘ������ߤH`��8�%�[>�2v��i�\��(���r�*����D4��݆1�ጬ&��	�ҭ����|��f SB��5ϯ�<=7%��8�rUa��ч����$u����V�n�����~cx�?M�;� �4�8��������}G�D�A&3o�So�l=4,����E�G���LU�x���;gr���v�� eN�œ�..�(7��"���G��i4���F�
ٶai�i���E9��b��S����m/������W6�A�[�V9/l9'�,�r����y�`vC]���8gX\�@V'��X�	�tb�5�5r���B"�z�s»���}����;�q��Kl!��jx;y  ߼R�8�W�Js����SIVp�7@�4�U����E;�<� ��v��u��AR��>}g
����n"!{Q�j��S�v-�ED/̉T��e�������}\�T��y��U������A�O�m��WPS��|n 	
�e�u���g�������eN=r�U!����[|�w�o�b䵑��Ѯ�_1k	B�{,,Qv����Ԟ�p]��V���gD�'j��[��|:�d:0��,�	J�㋟��=+5p2X�����L2��S����^��K�E�J	.���S�O �?`�/f�8	kR��o|-�%�I͔ż�68CN�s��0��*�cpB4�;Kl{j^�DE@�sЪ[n9ڋ9�������6JH�-�#x�ݛ#aC�a��e����#p�á_�N`�1ـ�H�k�$Τ��}4��}�G_��s:d�%R����|� b�mdr��P�JƐ6g��*�и(�8f�����Ȱ��4e�+s$�J��q���;%!_nu��'.A
�r�7�N��/��8��(/�OK�?	7�A���D'@���='�+?�Xn\׭��x]tk�cq�x*���dW���H�t��:c 	���2xx}���OS��Uȳ���Ϗ���6� _��;;�nE�ϩ�?M��M�#4���T�VܻK��v�%��d9`��KVZ�/�_鎿*B�dO�۫k�!�%��Ę!�i'�P�%_�+��F�%l�&mth�ҕL|3��w�ڻ�ۡ��-��}D�B�4���]�O�^���}<x)�]X5��[�+۰^���F�_oNŒ9��YS��_v8�.�t�3a^�PpWu��ȣ=Ձ �L�޾�ʱ{On��ir��u�]�	���CFZ��T�d��YijB�Y0$˓��,V �Db�$�V��/�mb�K+��r2�<�����T�k����e���ͿX5s�y����n^VI���1��2{�<5�/�@���m\�g���)6?:La���+�<��h9�E$ġTiX�M���F��2�ᤁürY��.�C/U��dX��v���*9|{�?�}���ٲ��}N��E�q�����,��P���f�Ձ�������A�;�sc��`8h���M1��m깝�dj��$����T]����2�����}x�B�a��`��"����t����`ԡ=����l(�K6��;����V؏]���<u��Ml�5U�7��OS�s����q(�[��J.Р P�΀��Ԡ¼%���2�k�J+���h��_5�>��J'� #�2z�A���_-�Y�`u�Ҧh5hK|xky�%�s�H��Ƿ�u}d���r�VM��$�ϯ�bM�hT��`p؅�>��w�����R9��r����f�Ǥ \����u���p��T,���#�a�"�,�_iQ+U:��#%
�_w��\�s�/��nh��� j��/���h��<�/V/��F�Ӗ[�����#b�~�	��o��jHP<�x���Uv��8�C�s���(QdA��R?�j'��<�"�k���іT��mk�}�ZC�5z��3�'�]ٳĂC��ӣ[��3>�Z��=6��(F��(�k��3� ��⢅%	+�Õ�11�8����44�A��ǃ�5��1��	�^x�^�~���u�w��|��\�qȩ҉έi�ܡI;d����!�ݟ�����:�n�G�NQ�1og��%�F���>��!ܦNBS��t�����Zh��e�/�;�]@�p�4�?�dG�O/�[3�
�c^��x�x!���Y���d5_�����8!��l�yA�ʽ=��9�I� ��l,~��h��\����p9��K�V�QW}���1D!�ʙ��Rب5�)�+,�	�;Y��������CPTI%f8�๬g��� �+J�pd����}��L�k�]ͷ�c��^ �T�����X�����5�x]{��2�j���l�'�A�P['��<�UJ��j���CC�y�V��)n|��]��4Ld	ˌ���'f�TA=�@[�[�c�=H��
S�&J*CsJ��t�Q,8�t&�T.�-N�����4�PSܘ��d����Q_�~uP���F[�A(����	a�~�4��{#�m��c�W�Y�@��V�+����;��(9[n:�;� |	��8�o/�Fm��D�����̠3���>������ ���qyԤ^[w`$�/׋���;�+hi�Gpc_�����՛\L"dI��H.G��\j�8�U�AՍ��ꥫ�ܱ����)ȽK������k��N:9eVw�o�=JFE���wb� ����Ѹ4�t����/���D2{�I�S�r�Z��^� F�7�%�a	I_�\��-ʹ~��t&�eY���L,���QoOcv@e:z9)I�(2�Q�5�F����ꐢMU��5G@�����s�d׺ny�E
m��t��u� �X����VOߗ�J�յ�L?���AL]�����\��%�i���X��4��`{;'4�H�ʹ�,���A�s��N �a�~��Ҹ�>f�Q��vo���Ʌ}m{^�s��Aa�o��j�0�mPeߔ�6�N��i�4%���%i�F�B�Դ����X){�Ym�C��}\_
��ћA3X��9�+� ��k��ub8���L�<�`�uG'�څJƚq.�"��k�������G�%+9k_ v���߿����xY��=�1b�.p�pA2�g�K�R����y�p���(�����ֺ5�'�S�w��H�rHs���q�8SK�4�����MmӨ�b�+,����آ�a���v��(J�K�n����CŖ����"�5��s_�uHmqu��]��`�~SN���wu�h�`�����F�;DX/#1��
1�akCV�:cx�Z�r*(J\�o����;+�.�;2�S��J�*e i�;;�c�#�K��̶���g�9�������u��;�y����su[��\"�x�a��!��̺G�YZ�U�X�C*��A .ϻ��;�w+�:&�����2����R�a�3t`�̆Go ���-�mqWڷq��g�z��y�{�="�Ƹ覯/��L忆�h.U�z�5�kw����:�: ǒ�'���O�x��Aa�$��V �r�ER#�'���S��L�3�%�()�rX�?6��u�bl,y��k����J-���U3Jn�~���v�,a
װ�*��6�Xl�IHoǓ �;!v�.c�[$�nlNIM�����������zu�T=l-�f^w��C�Րz�c4}��>��&�E�T����4oX�\#ь�Ol{ � �ܶ&�.L�Z�z�k2��Wl�.�Q��k ~s�X$s�U�p��k�b�LG��GV�0��⩱�)��k��a�.s}�g�h����ʣ��
��B)�2��m1_�,�<��Yo���<��Ja���Y�*=�sZ�pP9b�$Y��w�%�A�b���|;3��}w]�}��e�ȭo(�)�k���b����w�%�����RNC��8�������/s��P�|�iiI'��9�Z�v�pQ����2�0G��]̋����t�#�rW<���Un	1ܷ��yI��D}+rF�G��$ܿX1�r�z���*�������%�O����rQ��`a�fx�l���#bIu�-��9����e��xգ�]���. ��]����a�_g���c�(���P��ȯ따2�b���F�'����)	�����,5�+|�U��i�v<v�?^��3���Ȣ(1�'_8�^���\�<���
�}�J8zg1����t�Xz0�DD�C�Q��S�����7V
?�Έ��m�{[�~�;`�9U����`��_�lZW�h�_��!�΂�V�/1��E�/	�;q�v�(�2��8��Ti�kۙ�mK<�,Jd.����hKYa�-��=md�{��"uđb�7%Oװ�t:W��&�(�k��']A]��ȋ�g5�7�V؝���$����dXQZ ���\?;��@��=6Ѣ��Ŵ�����+B#��=��22��+����5��S��H\�[O��q{#�}O��&�n�]f2vE��I	#Nf��,��9K�JB\��DU��2�R@�ڑS�.I���B�}&כ��R�4(�/�;�kQa�%4�����s|��%�i�k"�O�����b�ۍj�⪏e2�vT�v����V㈏ú�<��^�E'E
�y4VP�d�>-�LzR�)U��,��\-�X��H�%Dҿ����T:yq�3Ȃ�R�Hv9�Af������$��h@2 �+Զ��XH̅FD��������*=ڼ����|��QJ���~1͕c��9����>8n��ג�}%5��d'���&�^]VI��J�j�W�EH�Ւ��HJ���R�?M��=�1���9q��XH�v���+���2,���CX�� 4;ݲ-+c+�\\�=�,}fI�z7�fGn'Ns�+�
(��$5NQ�6�� ��M�?3]�A#���}5J�f�d���YA��Ok@3��!J.��w�Z�e��Lu���3c��)+,��Q�P.��Lo,��X0�6y����m��wGzkiWIo�XU�o�[?C��n����)]�J��P��tR4��w��+!�&��1�������5��[H�H`
Z
i&��Y6 �1�' A����OAj)�FD]�4��qT�aՅ0�{޴�V��>�w�� ld
<-H�E��-2�.+�dM3��)�'��3�
�p���?��B���ڞ����:Yh"z��L�R�� ƿ�Շ���=���wb2�ڒsѷ�T/M�����&������i���և��	�FX���t�����
�wۘ>>�5.�ޔ3�y�߽�m�[5N��D^)���q�N���Vi�J�rٖ/��(QW�x~V"|���$����DS�E�5L�I����[R�Կ
�����f% �z��7��A�֪��@��U9�z�v��ݻ)p稶�H�ei�䨰�uSm8�8I�n�̞N7/.sd&�4�:��]#�j�su���~�J�.�hT�S�+$��mԅ{�Jtpʹ*h���r�^0�GO�E���5��/.��|�x��9�y/Z��Y��{�@fG��#�v@؉)����0�lDfU�dt#�M��D���^B`�,��;����ԙ��_�l% V��l�bX����M(���}���R��g?&�Ss�qr�����gXv,!�$�:�~
C���}ϲ�C��g0�o�����8&r.��DѸ������o�[}�Q���yw�	�"4D&]9mc!�ʵ��{�';	H^3�׫�d66��D���U@f�{g2�T'Ci���R�-��y��3|�߾���>EՏ-z�ȋ��0y��ޟ����-a#�C+'�L��+u3zp�@,m��j��{)nuW�M�j��z�)�(��Ⱦ�����ޓ��4)�.�|1�i���`a���<2X28뷔�%�t*�c���	�����X����g+��W%���1\)��C+\6ATG�I�5�L�g�^�K��N���`��j"����uS�`���~�~�e��R\ϻ������&/%A��BZ	Y9�T����2�"ȅ�K®�4�]�1����b|��;Ec��ͥ?*u���5� ��&��#
�ҹ��i�k_�0MB�΋�{�u�h�Qrz��M��q\J����d|�����=�dq����,d'��d�2����"�������� �ć	��篛3��>r�6FZ�yi�z)�:�CV���Qabe��8� Ѹ��� �SA�(B�k��eC�(�9w�`��DE�%�'��E�1�q)�՗�Ǝe�������L����f�d)sMg����Z��1��Wz�����^�C�'��:�U
Q�����M��B�@q+Bq�s"O���.R!?]�P&��~\�}���Èb�����r׀<�z��r�]�K�4I�IC;�)9jU*�ِU/�Y������]M��Ó�q�i�;����׷��ur)6���A-��&s����Ms�d^ڰo��ѱL��l���M�DA'���7K��6�h���T��u1�X�þw�ئ�����p���2�x/�+�^�XM��S��À�l\����*IR�������kՒo���2�/�ӵ�����&�*�<"h �V�� ���Я�H�o�&<~����(�<�B���3`:�͑G��7�Z��S=D8'���SΟaP�7�@c�0�r�K��	����Mx'&�H�a��6�v;�c�rN���B)���nE�i����&Dw��,
�)�:���軅{������o��j�.%I��RH9'b��0W�)��W����G�����B��6{Ft[�~����rez��ХϠo>S�-�!y�T`Z����d�٢���_sÄ�d^E��������>-�����������	F���4C��֗w"_�cu����9���c^�վ�?0P���1�ؾ;�m;��DaryTa�a�F�)D�w�ބ}JY��݌��G��KN�E��ԛ\vv�2��'���Ǔ�-|J���IE�	�[b�X���ڻ$�Lȇ��]�uȢ�CL�M}ԥi�����3�[Z�b�˫�VO
Y*�p�0'r�" �O��7�S\�pC�8�>����.%NGXF���>s.keq,�b'+��Z�gqg�y��}٨p��\s�|"נ��<�� ����������6RG0Y	a���!�'�^�6�C�����V�.�yS�.p^�,y��(�����N�[2�\�ӂ����|���x�*I���o�b/�e�u��"�����r�;J,]��1/�������E���d�k�q�]�W��}ޒ-1����m�XѾ����^_iv���?�������*<�h��?�e�M�����!E�~�X�Ç�ճ>v�4�=h�X���Z�JR�{J{�R����;@�H�N����o���͂�
X�F9�����(�"To��7��>5�5[��ޅ�7䁜h&�~'�|��+�G>��h�>/o":wj��%��D�M�yM�Ha<�T�V6���
��YŬl�|{�=��K�b�ja�ҡ,�� "݀�p����/����6������惡����W	�����|O�J�D�1��[L���;?y��Hy�K{�[������@RF��+���gMr�_�4�U�
�V��!n	/��ȫ�����zR*g��hG����iΆ}�+��x8˧%݌u�0�zeZ��+ B�\�'b4D�i�ۛ��8$����^�d��?����ahI�F GF&/���r��i#�{~�w�y�Ǿ1���li)*�ҫ��c��`� �Ҧ�y���^���BKe���*��G��f
 �I(m�OLSWL�u��0H���z�}mW��ɬ�[]��ʑmZ1gWw�̩<OX��X�0Ae�AlѠ�F�{�m����B���>s��������� �;�R�d��8l>hi5mڈ̢
�����2p��c�&��)�(Aӕ!�6�_&Y�̙�	=�KG�n
�=�ެH&�$h*���yr�j* gș��{��7����;�L�~�-��4�W��;7��pƆ��}�FL�35dD�?c�\b�nq��f(P��;8�Q��X�J�����Mˊ�ej$�̢���$�~Qǝ�`�SUWڹ�f<�`��S����z�
�Kb�1�n6*?d��F�d�o�S�%G�5�&��1�N����U�[����'�zӈXc�1:"9��,0G['���H<*�'Eh�@�*�?M�.�n� �� ���g�E�,�J��a����+��Z���6���	m�2>/�e�hƌu_YQ9S�WuC�}ɖ2K�[HJf���l�Tm9��5�~�<�el������Uc�9�e�9I���3PG$�5#��=�S�<��e&,�����7�"�t��4�,o\I��i�U1���/¯��g��Hޘ���O<������!�_g���jp�Ԗ����,�w�7J�7�� ���֙c��)�w�Oo�z��>ڝ��_�U�&].]G��{Κ3��"�Z�H�xk���gj�S��!f^����T�䍏�Z�.{����`�fC�m���S����0 -1�D�N�Q���p�p�"��c���x��<�0�����
D_?u8�0�<|��
�	 ���郉@��WD�j�y�a�r���\0xn�����C�*�վB$0���J���u�8��}�D�:0�����9�����������cx����Z�>=k��?P�F���`)�������W��+|���͐!���/�tT���E�ާ�E�!�T��;��vח�dK���տ�q��Ȼ��{][\>lیg*9	jW�mK�2&��y_�q�Ɖ��OA�ߠ-�8ٙܫ��ٔ
Q����\�L�!r4f>D5<�<�>��A�rW˧{U�JE�ĺ�3�AF�F��@���i1�%o��u��;E+d@���<��p���XӚW�ǽ�2�UJk.�X��o�hY��"�S����u� Os� �M�_��@�n��g��y��
 99*�V4d̎�����O)��р�:��"��f!���\������XHx���ڦ6L&[�g.B�I�C\.�Jjx��=R�y��]i%#Q4צT����?ĵ���,��H6�$Ri�0Sja~g~E}��SH��hH�oF��� ����*g7?�+̽W	��uE2M����ޕk�8�)ij����a3�PX���Q�|o��Vx�M�D�m�����'��ͻ�pfy6�=�
c������#v��M�[�$)1y9����HK��UQ�F��<��J�v��l@u`�(R�u�5e�%�<
֏������B宐Ƒ���Ӱ����^C���S�S�RH��Fg�bIv�����J�	Ʌ����2��3l��� ����R6��-u5�bV�Q�&��PsP��DA�Y������jJCq@�7)��)nF.7K@5��(�e��v�z�7�l!��I�|Pʭ�u
�hܻ�*�=C�F�}���S�ŅM�/5AM��U&������:=W���fꗅ���¥Wt��C5���G�2�(��u0Y���HW�4��9T�:)�����ck���jj�`�5����m3C3A�2���iPM6��k<He}�#�wH��L��K�	߃m��s;�������k9��ji]wx�BR�םS�<�,o��q �{�o]Ip	ڳ,z��SI�_�_�R���ƑG%�SL�T���������߃@
�g�ԦcD�V����j�j~k^����C���+٭,�"�epS��'�c��{���W��k*�Q��ׂ��zYHl�}3������lv��
�b�&!��Е�8�{��4�U��^�,�	�J=�h�6RBK	E�~y�f_7��&��\w�"��R����2"4������O���Mi�&D���~���1�8�ߚ���]$ȅ>�`&��;�>nҦ���C�vw�G֪2n0�~�[��H�^�F�]
x� ��h�Y9�'��Q�@dF~/�+�ؒ�h�v k0 �7�	4�4R��z	��_Ρ�@PUM\Ͻ�4��
��odR�ZE�&5���o*+�5d'U��ƌ\��>���x����������Uw	����=f���%a����kՍ��=�q�dc>#7��K)���ڬ3�B��Z��`A�����}ҳ�c/!D@�#F�6�횓�;�TK����|c>�ed���y:BA���n�����qDeĝ�j*#uN��|T0���"��)$4�yGyLVG9ѷ�N�Д>6�AL���2L�8�7�9��q�K|�!�kf;�n��=���c�V���_'��C6��vށT���\H������R�t��.��u�E�I��L�}�̹��m��g-? �,C$;f��đ3��A$|A쁘�~o�i��8��Է>q���7W<G(u�&�1=�&Lݷs��-�������T �խ��V��a (���,�<�o%F����䣎-��/�\�]�U΁9uc�x55F�x����{�EY�M]y�Z0���ߺZc�����z�h�H�ɿ8����X~��T3Ka��z���#�l6��b� ^3��7f��B��jR
��:$KD�؋��AA���-ЇRO��/}w��ǝC�zV�_�'h/w(n���6t�3^;P{�����m�m����~#~"
�
������I��ܛN0��l��tU�w�נ�V�y>
 �\	On|qQڻ����	ƍ��n-$ۍF�/_K!��f�0s�ߩ�����4��4Lf���F6ĭ~yv��Q3���QW��Tv嫯{�j�^v��`Ɣ��`&��r6E}c�ƫ���C�ܾ�p���UV�����M�g�ڟZ?MO��"�ȄN[���z� �����q῅�FFH�)0�5����\?�-_l�,���ŝןs"�u��� �B($�b��&��d�Z$G��Q��r����
�M3Qk��(Z��$�|��KR���1�m�>IY?�i�a���#�Y��B�SA���Q�{-fu��=r�k�R���2��R���	op�T�F�$�kw�,�{�\�h��Ư��R��W�����6��1�;�'��#7z�&�xA���N|����DT����1����lt9�I��>����3WgY�5�S���wK�D���������J�[���a݀��'�W}[�/�Cb<��	*�P|+�BW~<����~~����Y�
�Ǫ�f,�ZD����_��,�ޜ��/��{- �ƒB�~ZU%�.Z0���!-ejX8;i��vu�$��YS��Q�|�E'n�!���|૛��Y"��ީ"��}�Պ�+��P9� ��q��砑H� ��a�#���`x�KH�Ϯ	e!�x-�*B��n��~o �~�3ڍ��X�/�L����*�v�YTo"w���7OL��L�66�v��1�I�����LAC��U�儗>5��剛}�7�s���c��vCI����)��U㎋T�𠅖�ل�*'��s��8��Ք3�����K�ٴ�<$��A�.]�f��-\TvԳ��҉V��x)B��d�*������~5�|"��r�h�L��}rG��O��"$�zV��8n��:�;7ՓGYæ��V���$�dq�}����w8��L*ν�)�"IΣi���a4VQ�ibZ��F�f��{U"�a��poԧf�F`��f�ş�Q�w,Q�1����<8�ógq����!0
}�r���G�/_�]X�ؤ�ڵ��cecG )	Z6�d�	�;LIS���jl�ɷ�h��V@�m�����L�O���eO���◫��P� ��l�跩G�L炧�Y���>}��m��:8��0r;h�\K[#�B����P&�����f��R�uz�g8�%��s:�2*�JT�?ݯ�N��
��J�M8�k*?�]8�Ԇ�1'�6+x�*S�	���s:wB ���w��XL���4@o�ݍ%ʑ)��t�V�M���,�H�o��{[|W2����]��̕��9ҡ��b"wl�.��E����=L-j�rx	1��nK`M�����L# ��]k�� ����V+[r��"D�l=a��zC��9�Cuj,Cq�^��=��w��pL�� 8*�N�cp��uD�r���7� r�b��+����ь9�Y���o��5|";��X��L����{� �bak
Rh(�|n�E<���;�;��#�T���E�3�����wX�^%��
��hЌ�ud�� ��c��p�s�^�[0�9V��EI����E-gL|hA�t!*��.��Ъ�	�u|<m��`��!��Ol�����8!�.>�l��]ۧ��ʭ��@8�t�uo�r�+΃>;�׏`y�ƹ-��OL`�S�i�L�Z`�c�?̱Y����B��n���d�_5q��Y~���"��Dp�����	y��P����m�K춆0u��9�
�������ϛe+�>,���w$�b�*��EΩ��B�s_c��G\�1�G��iB��c 1��GQ�j��3�&��+W�G��%	��'�(�LshZ6}G���O���۾��i�+~W6��[}��fD��̡�M�=x�
�ߟ�l�q	 ���Bh A�y�+ϡiB�5z6A�վ�"84F0d�5��`a�x$ğ�C��ޱ�f��M�-�?��F��T:/Ɠ����!�I��wv�+VW���0_P�" ֚���(�ŐK�Lcq%G"~�`Ol��˺���F��Ҝ�<�<�X��D��y7��p���?OB<1��i�,,W��T��1I�t������&��W������?%�4��E������@.-}~�����\�����w�����ڊ�)��J3�vAp3-k��{�AJ�������6�ww-�u���r(�3���}�>�Jk� 0��qB��bX �椇����Y��� ��*ue
p_eBGR�H���k0w�I�q}����6�kb�C/��@ط����V�(d�����tG`ks�}�X5/��8�m����J�ߤ6X�����ߩV��䞹pˢg[���<�ˉ�Y����g�f��
�9۟�_��! ���q"qu�X7T���0Z���#�U7�5+��p�ӾXncl��*�vM�ˍ�@��$��b����{T����'�A�?S��KY7����E}͖DN<�7{�������{Lj���M��^�$KD04�����D���<��W%nk�N0�^k4f!�K�0J�6�l����1��~�Ƭ� $���O,C?,vB�2s��4�OPѧǎ�u�*�C�-�,�#�D����7���Ҹj����u��)��3TG;�����:9N�����Hո|Z��7WbHI���>5�+m��2�{�g@������ڻ��_����t��f���F��̄!Pt[�W���,�hj�CV��w}��o��k}m�b����s7u�yڐ�-��<rl��^U�����Gb� L�[l��]�(5�m�7�`B?���"*�Nӊ�.����,:p��r8xKc�7�Ҁ���dÛ4�Bx��� 4W�E�"��lV^�F����j�Z�_%���қ[�Oջdj�!l��,�}Wn�H��s�8|6]G�H��� ��+p��nJ�z�,�\=հ�E01b��r�C�|�����,y
��NL>ۉ��@*�Ks��-��Mh��umd��0V����v>�)�w\.Y�-�P�
f�,W�ă���� n�M?����8KD0�@�%�D.kJ��$~2U'+��V�:��U�M���w�!ͫ��v��=|&/����\�N6߄�%\�1�>k%I�a�R�����^}�2�#��n�@L���<�٭����j�ָ���
_�DrL���t�c3�=�q��!�_W���e 7x�/��Z:�'#�b��.��a(G�aN���'w������Y�
�CMs����eƘ�
w,�,�>�T�[��Ќ��=0�!��0����h�`�(���h�^��w<9Sv�%�҄~b��rL��L�~���z��%B�������_Ǧ�\y�7�����M[��\'��k���Ji��튿|���Nx�mk��>Y�/��{���xj��Q�k�Ka^�!V�/Ò-4�c$� S[�պ�C���
����}�U�zk�.���1X��G�~3#���J��.�#�U؏�@�x��ZҞI��&5����L��������ËY6�'T��x�Ը�9B+1�j�"g(Lb*ܨ�xm�V�A�n��d]���{8;1Y8��ds6�=t&Փ�2@9�X�k�X@�`�`za]I�������=�uE�p�>GdbA[B߳���+E��G�,�p���<!]��<���]�{	)�¿�a���������eq�&	(���L�
]�ʕ������v��.=:pa�57��z&�{ͺ)C��~U,��e�< ���-�;�`�w�Z�t辙ImBI��-tdECK��΅�����3νB39�\����ac{ղ�|ʦ:Ȧ����`3�z���_��
#m�Օ����6qU�Y���.h�/�{ʤZ%��	{U��PXx�.&v%���b,��o=!?��ޟ�����F��EͣD,��1��!zq��3�Wi�A�Қ;v���ڛ��T����2лC�����![&��̧O��`t�5��d�41��L�ȳ�s��p������?�g���|왣����B �	-�N�!k��,�υ�y@�4�}kb'�כ�`ǮJ��̡�v ���������
d2M93qR�ۏr��v�����$X���Ӷ	p���n?�+�[�Sd��9��
iH��7,q�4����_z	��P��p%�j�y�z�­�h����^ޱ�V|^;:6��C���<e���y3�Y��J#Fx��ʛ��f>��F��<��Q�t�އ�����Uu��P�����a�J`�gf9 �ڧTqѭr�ow҂t����.��&,�׎��м�#[9�X��U��,�K��fT�%�j�p���F}��.a���N��~�?���yɠ�-���Df<$ʴ��ԋ����� hz5,����yz@�&s�����3'y4[Fw�Ve=Q�HW���e��9|ۀ�YX���md�
����f�3���Kq�~��U�\���<x^-�<�ҡ��q�0�K-A�7�נ ��y�5#��<~Gg���MX�ߞfb��!���y)�1��N_EA��o#�e����r:DD,���B���]�ZD�۔*���ܠn��&u^>�SWH���gR�M���I�^aCQ-�B;.�'�,gS���J��J��:�����s���B޲����W~Ck�a@\F��=td�BQ.$7;I%~m���}I()�ù�[�x��Ϟx���R����	��n���Is��g�(xQѩV~i����y�mWQ����O)�� ~W�a�X���W�*�dt���Ĕ���i2��]E?�/=b�糽�Վ7�JY���{
�ڤ*[_�;d9�����A��qc�D�0�6�G��M_ht1;�Ԗ�ln*G��6�������F���G�<Y�\S�Pz�Pw4�\�� 7�X����b���>#e��ci^h������]�y�m�.y/��mZ�p�m�4l]���tˉ?F�&9�P�d_��7͉7��e�ଢ଼QC-�v-kp>��ᆣ�g��akc����LL\�j�V��z������TW��~����,d����*T���ON����������g��	̘}e|�b�q��pm :�;~W�L/Hl�09+�^�-��e�lZ1Ȼ��/]�J�1:��%�b��e�!0�,��N�Ĳ��X��y�g�?�C�C��O/j|�T�P��m���>{$��ř#'E����Tx�-芙�饐B�lȼ�I�߂M\ ��8��2_���Ց,f������)�@I&���;�d�GC��;��g�YxT����ӣ�ȸ�5n#u����i�O��mȿ�AU��I�g�A��j]6ɜ:P��C�@�I���Q��h�D�L��fY{J:����8&����Z!�V�h"D:S�����
0�Mq�03wd��x�}Ő���+�s|7�|��h��1c�K׶b��ʇ*�$�-��9����
��E����T��7q�]�(ʺ�f��h���x�
���G��8��k�7��fjr_�:nZ��`����Ւ�'Ǆ����>�a�m޻%�W�hV���GbiV�C�B�n#i�آl�Iqr+�y�9l�M�I��Yk%o�ɮ�"�$��dONM�#����W�']T��J�	�"}�'Q>u���B7n����6wWT~ �8#�C�u�KJ��i)�	�C���$d�D؝��K�c�P0��T���]u6x���F{���j#$h؋���_��{��L�y����)��IWUP�YJ�<��e枎ӡ�5o��o��Esv;u@�#G	��0�vie�%�m�G�in�ϕJ'bh�Xv�G���Ie�������Gw��2ž��t�����u_M�וy��<>�����L�x���d?Q��<���J9��Ɗi�W?��ȇс���l�����8���wߺ{�-�'l�.CQ�n�ﶫE�Z����5;2��"��fQ���]O���'�� ��lM;���+t���c"w;�Z�o	���N�Y*�Wc6���C�?�tզrg�_R�=Y�Chb"ϡ՟ֿ��7wI��x�D+�!J[k[X΍��E Aс�LC�ib���k��#�g��`$X"6R�v��.�ݜ��G�˝��.�y�5թ�����}0�p�|�	∧��E��t�/,5`P��БsE6���[%ʈ��O����d0�_f2Ɲk��+� и��j-,�r�3�'�kb�3;�`k~���B�!VX.Eg����@�/���"���hxL���i`+��pp�ٙ�\$��`�!a�^��Ǹ4`K|
�z{-`������*.�S�d2�����<D�����A���/_��2W�f�e'���8D%��9�`M��8X�ְ���2x�旹Mb<|�*Zʄ:�����	 B啁x����P�g�����ڷ��"�#XY�Y�y,��!S�9��E��'�o`q^���Cү��6�PjB�-5�+y0����L����)=؊�fH/�(m���GK�����'D`C��J=���܈�y˫ᎉ��P�vW<F:mjo�$�S,��]�"أ�} eo0�iT�՜L����I/���3�L��T�X,�XX��!o=l���X��/ZG�.��iU�y�W��Q��q[����������[�.<yN��{�1�	��%�~v�l��T�w�1M�{ڙ�	��m7ȻL�A������O'ђ�m	L���(Q�`3��Vü�{��.2���s�����5Y�|��$G�$B�G�6�%�z�ǥb����5|C�%�*J}̱w��!��Gq�z�	����q",C5���{����]��4mb�Fi��=B��<�9��U�~-���rb@ql$�<�距��?#�.�Sy*;.�L��p��ɲ�Z��|F^b�Q��΀��%���t�,y�oCc�RZV>֙i����t�.��O%|�}�|�fw�C:zP��$��Q�֪0-)��� �Ӳ{7C�lwViP�?�����D:e\r"�
�����v��Z�P�gk5���2��c�͸.R�̅!F���\;�X|�P�.�jj	�ȹ��Ū-��}���bj��Ғ���,�c�-z����E9* �j�K�0
˟]ɐ'~n�{���#Ց�gl�L�J���g>l^�Y��d�%�&;܂�aD�b}��?�
�@��C���&�@䭺����&�ѷCU!p����"l���ԋ	�����P�b��1���#����e��Ը�p��a%"�û���n
�y�3@`�L��2�$-)��kh�d�*��4�qP ��]�Exӗ�]���G'� ��V~���[�B-]7�͇��:�ž]�AʊX���'�ޣ�c�S�}�y�,�H3�шz�^��0�A��{���ضR��<�����W�8��<��D0F���n�gI��hl��<�`י�8�a�����@!����� ��M$X�|��Q�H�<�kS>�:���A����9,������,JT��ֵ㦋�ܕ����za�Z��(D�N1�'��)=��l���r_�_�~��O�XS��(@4qiFQ��Ԣ��5�l��vL���o��������D��Y!-�hKF0�Y�X}�+[��-�``��ׇƿ�0���V���]�8�jF$E����r�[�n���Y?o�iF��%�$����*�5�>�Zp�f`���?����p2;��5� @`hJ���,l�ٿ	����(��dy��|qgi�^��j��!UX2Y6�t��pX�/�R^
�<�G������Ǯ!qf���;��5�N;�ʔ��|ہ�uyQ_�Ԯ�4�����������W�h>L��SMvHc�����D����J��M��N���A�
�Rbʨϰ��3/ 7�n���īn<��@~��f����.Y�Qc�����ˮ��R�%�2��~.g1R��B���s���̀ƣ�(h��Z��'Y0�0���{O���g����ϻI���p�x�KQ�?���@^
�i���#���<�S�_�B�Z��V̊�.$(V#�����}#�:*�R� ( ѤjCR0�w�K���5�6Gx�C�����Ҥ�T��+2ΎY~����	��jW���@�Vng"bJ%��¶#Ҹᥦ�
B�� q ���.>,Uo��(o��_�n�,!ͥ���\�$��@��z��VKT�����-5��j�?���]����]�������0���..�n���S��]��GTO�~VM6���ȗJW3 w��W��Cm�����^�t˨uٜp�xIYl����'q���~�*Nr ��b~�r��S�DT=�&���PU�y�5�L��z�|� c��~��<�=���^c:��ɡ�Z]'^Y��<zE�y0��̒3T��m�����bݞ�`���\S�)��\_b�NO�}Z����W�O�������H���wh�����!�S�e�ȒO��[�b������g�9��hԭva1+?�p��o�������&{ޫ<[KY�D_�,ёa7?}��0UC$�L�cץ�M �x����iFI�(%g:OӖbFo1��3�^|���q�u�"\.�m�K�G&s��
ww �Kڗ���3k]V���z�|{'�!,���aﻼ�p2�}��Y��'pI��v/t���r�2�X�J�	��(�2���r�����Y�~X�d�~6G�)\$݀�m�?��B��l*d�F�W;HRW��^�DFUy�����>"l�Mݥ��L�ky���`��	h�uj�h�Xȳ`�s�=իŏh}�IU���S��ν��Ӓ����V���=L_���M��!�LU��:��/P���Ԭ�L��/[M,���#�y�_��5p�5��lg)Bu�M~j�=}����d�̫�����6'Z�i�Wo��di�J�)H�{l�rK�%�p�̩�uw���)4�d
���P15B��P�[h�Ng~������{�I,�Z6�Eu�=���H�`�`���eXfG|�h>���Z�Y�k&�a)�_���H̺>6�g�g�W�����D}���Ĭ1i�F����SHBX�69S�W�� ����)��YRS|�`ņ�&���n��W���KȖ�6lYt� ������E(܎�P��|ޒ�X������V@I�y�U�+��C��<M��A����R���x/R�_�����E5�>~���f'��C2/4;S�z�$1�5��6K����~.[#=� �`N����!x1�h�kj�qᙂ�xU��K�\����!E��:e"f!Ow�rP>t=�6�yf�6�k*�X��5���o  �Ʊj� |�]�!�"��SJ�U�d�� U����Ұ����x���:%�ys��y�Z��@�.0�u@H&�6���� ك3�*{��ƣjVr��Ks�sXE+���۾�+�����4��3m�ȇ8�C:[������oN[��;m;���H{.��;]!�KVS�����$?W�������Q�S�y�hǄ;�'��'�b�w�h����[p��Ƚ�<��W-��^�D����۲�3ɶ)yu8�y�Cry���aL#���^}��|�y-B�[
�ś�D2}���`�YW�t񥀷��.��q
=� ���Q��(�f
��T��>�/v3U�3�<���f�yU���׻��@�\��xJW���e���HN�%�r�7������5w��$��9U���.[���1��u����E��nn�����������X���'>�%�Uq���E�*db�O�ۻp�Gg��n�5f'bMm:�O�?��Z�	'����;":�`���9'��:5����Ky�� ak3n%J�k��o�]>�ie�)y�^ ��`�z�i�y��d�a�=ǡ���(99���1i^'k?���H�R��"Y��g���Mnb�`	J��G���lî����ڙ��6�P�ʇgG�^n0D��#f�)���F�35+� �l3	L�.�JF�%*O�,D')��u-�B��2u�}<-x2��R<�@:��_`����F$�w��T�A���Ef*`�bY�5�|E������?Z*<�LGV��˙H��M���w��n+^�J�J��5�P�$>�##l�O)�t,���[�>I�ݖ�=�1y�4>(�e��_i��R}\AK�z��k��0փ�Mğ��Qr�/���.i�T	�^q�<?痥/���&�s+�g�.����s1�[4I�)cUz��]RM������;�CiZj�b�V��׈����� �Wf���B6.���\!���x0�^��M�+8|�<����R��kV&�]ZY(}�(����m�}e�q�q�sk�f��.8�&|�O�B��c�Ms��U��������k%W�F麪�C,M���"HF�����Ix��eE��!d��7���A/\~���z(-�kkR�������9�,��_�9;��U�`�$��7(���&���笲!z�,έ?�l#KJ7�hh("nx��+���4�����"�Lֻ�:�(k�@���Cz��z٫e���[�
�t�W?�=�ؼ�I��E+H���$پx)eM�c١��?S������p�Z���ڜ��$�h�&�r��I˙�8�cu��ڙ2aٔ=F]���R�f3ҭL����T�7�}�u�:��{���Ƒ�-��͇�]�8�
6�����E2�4�|Z[Jl�g�E�rN�!6�ʉy��m6Cyc.{p���`J�F���8mY�g%F�: (�|34��u�7�ܒ�c���"�zkC�Q7��˧X�O��x����$j�![�m��Ħ�*��O@�k��Ȳ~�/D�zn(���T��9�2�)A>�����f@D��e͵;k���q��IG/8�s����/n��+�>����]�d��� ���:��C��G��?����u��X@�a_��	��MO��pšo�� ��
�ɒ�{n��B��>�6i���zK�� dJ8��i����h��[-;��@�q���g������l�ڨgp{D��)E��DTPw�N	q��yn;l_}�ԣG9�&m�28fh��}�F�/Mͼ7�T҇�iE��Y����Y��C��]�K���(a�N��1�"�^8�up-5)m���M$%�������=|NT��
�h�y�k�z�,G�p�U�B�Q4Ѐ���I��� P��Ǣu�����X�� }L�����Y�h�����L=�)K0==eo��S� 2l�����%�����j��z<D��f��c�p�h�}���a�n��DU�K,�1{��ݲ�s�Ip6W�2�SȐ����G�	����r���nUeOC�̟٤���C[`�J����z��˰��G�=��A!"Ë�RuCf�0;��b���:. ut�y�� =�0T�ρ���$�L��3J�	t!�/�~1k�҆��j�/��E�F��}�<�ڦj{��a^�/�o��rX+L��L��͞���e�RX\����Z��G�.�:$��&9Fؚ�҃���n�Ԟ#�0�4���= ���*^e֍#���2�,J$��G��2��sF�_@�A��,����I�R����TK���2�n�/|�T��A�iǎŠ�
�MYIζ=p��T�
�i�<gsI`����11�Ə���׭���ޔV}�]<e
��篗�������8��<T�9Q����d��W^V��w	��?���j�� �7ʠ��0T% �����(t���s��x�[�p Z�%�Z?��Hswp	Y�SК��]�2I�$m �|H�k���&pΖ����A�]3�։�1��[���B���Q����Yjj6����֮�n:c�p,��&`z3����*�zԲC����~��\�[U�M��m�t`��
��VJ�0�7������>H�"��7��H�
�k���I�!�$]���j�����PW2㰢8�6�"b1���jC�@����W}�l������;��G���`R�-�$����?�Sf�����ϠY���������h�%�Z�S�q�ocH��A�s�È������x����S�jsa��A�eZ�h�߉H�"�Y4�K�j�n�G��j�9ܳ�2��Wm؂$������Y}!�jY I+�h����04Zb��z�X]�����x1i��-d�}���q�`�y�8�;����W=7N�(���ɦB����~\�v0�W0N��<�Q��Jv�q��4�ۖU��b�f��Se��jL��jr4��2�["���R��mv}ZW�(��"�tϽ��E�i��״!��rZ���_�����|9���#��HО�T/#��(a�S��-9k& ����>Z�~��N�m~��v6z6n�m�H����~L|Ƙ�ΉMa�`!�(��F;��?�������`��v�*�_׆���Ϝ��j�����!�q�%�/��y�Dts��DV�wĿ�DhQp�����謏	���ݩ��W�B��j���W�V���DSk�l8&(4�{������C9C`P��
ַ�N�u��[-��￝�^�����E��#t�����?�b��nց�P#�����z#�d�KKj��T�c06}K=�j��T����s�Y)P�1�0i�ϙ��|�!xf~���~�w���e�Z��ѯ��/����^�^G���`F��"Y\!k�&q�MO�e�ϟJ}��I�J[-�f����Bbu�檌(�x��6�:;e���G@�:6�Y���'ʖ��V���W2�����7�iW8��ŨR������%����BȒ;��U��)��qN�y��,�.�(�/&�������5e�a4;�^�rn2�v#\8T�D�]-��ɉ��&�6F�PQ2D`�M���R4������\W��0oi�Em���/+��9~(�a�uF��:>_���s�B6uy��I$��-�J� �ae�uMv��<��9���T�
~\���]?5�$�xkz����[Wi69WdS���]q{�y��%��vCw��N�z3�$�=��$�ն�ْ�4ʁ�����e|���L�C�{�_$	��Q>��-"��D/�r>;JQ�8	Pzb�]�L�Ol�ͺ����?0�6pr��h�V�/ȡ�<���c+jR�	NQ�_�����R���HǷ06��f>��:#��L�@���ڒ�d�qok���ҙ�N��Q@�<�����A������,��q��מ*��{���m�s^?�!WU	�b~��;���qyY��ǒLaG���$�E�%'k0pE3���K���0@��
��M.��98�&7�Ozq��YR=����g/�N���@,@���>�Y�î�!�NS艜���=�6�­^G�-q�p��'���]4���a�k�6��*��/�[���>�Ω?@_k�U��K���$�����ZeI���ߋ�)Bω���U�PF��xw�
;�.;;�t�ڙ�O۠���c'�y��s�Q+1�5*cCŜ�:Ͷ-����Au`%�;����Nq�z�ꖤ�y���o���Hh�����DO/R,h�l���y
�i<�A��_ŭ	��a��/979x�B3V�t�Hg���������S���ȼ�U-��kn.��i�JC���q;�k�i��]���<��y~���i1��oM��F&�&A�a1j�~�!h���D1Ú8�a��͂��FQC�W�:)l>��`E�h�^)z2�Q��jn�Y[�6�B7ú�9�%��b8���X��B���xE\�)�.�E��V�6����W�ɗ�-.x�6L���	��1�b|")O==�MO!`E�<�u��D�'i��K(lhP�QL[�{�Ś�.�|�qd[�Q�S�Хն�l������|7��+�}���OV.P��tK�'U�I��y$?*(��A]35�N�~�� �	�������m���I���0LXM:����&�K�H
��G�B,��ŏ~����2 ~L�3ޫW,:u45�ԅpnT9g샍:{�a^���C�R���B��B
������������5�#�8b.�?JA(��0�;��8�9`���\p]���W�loq�d�ٽ͜�\�W§E�rs��rz�ݡ���~�ЈoG�����z	_IWW� 4|�gͻ�x"�%.M6�Ud*�pU�F��t|9۹�h��2�o�K#�IPX�+����0����Z��3ɽ�'S1�$Yf��[��/�HnV"�)�����vd���z�K����]~�E���w�l���rx��2�_��ޡ��Nѧ���L �$1������gt�* oHV����6�p�S��:�����D�(pǄڝ�����m�z�/�v��XOk+�m�P�.��cN�} Lb��:�ܘ�t���Tu�ڌqDQئ5ل�rU������)�^52=����w���A��k�Յ������O��Nq�ra7�S��0%��p���{��A�c_���z?��a����-`M!�"s���m�fnTq!�Dǉ�u8���noP�ʃ��5,8�/{	���R�W��))A❄�����3�y��,#zޱ���\��0;��:�j�Vswv?%%�oW�����q`�����^<�����b����C�{��|�C[;��t{�S5��|(x1
�g�&����-��=��)S���W���,Nė�Պd<�3�����X�o>D;�k���;
�֨gZ2�q����^���>�`P	t�W�8�������L�-4O �3̩i;"i�K�B��QF���JϦh�H@W?� ��i]%=Pcܨ������+�0�a%�Zq��+P��Βaq5X1P�AP)׬Y�Lr�7fF�U:֍���HP����d��Z�.�E��俦�]��P:8�rq�I/ޞ2�F�;��]e��v��ۙIݐ�j�#`�<�^G^��C/E{����)ǐ�S�Y�O�X 	v�1H����V�\���B�G�mrXhS�����ɷ���:��yI"K�h�OMƫn�S D�~����(_÷��8�!�E��M1�h��Z�5�R{"���2���fYګ���K_j����B��
��!�M�7ۉ�j�R]
��f�zC腼Dü�������@�� F�����"��WA��L�3�G��L��9�?u;è�Y[�n͢����c�f�;a���7-?C�q�L��l�c��d랠YA��X��Aj�������~����5�	�i�[}?���*��!������I�IV*Όh/�GFj�oxX�vy����V�"�¬��uO��Æ5f���~���J�a�w�<����7l�_�sRM|1��8-��i:P����Fև�������3����9�0��
����վ4��sڹrd�z�2�gw���4���fu�v�
���p��'�xOu��]+�|w�cq�t��J�3q�k&rֹ����Z��p0�٣�(R�q�)v��=��T��9bF?z7��ʷ�y�۷����T�:	,V`�L�u�D��2j�Gy�K��v.�d�\B���|Y'� ���%�\���
�]��^&S"dFnG��T�{߆V�	���� �3Xq��٭ͭ?4�.�=��{X,�5L���Z���V�FE޶�>pg�0rfT��S��c��C�?w���_W���ٽ�A? �O�ͣ6����S.�������7{3���a��|�P��d�����58����#.�g�v�[��C�Vq3֔��9�^"y8���n�l��̢�2^��8�
1������IW�v��-�\v�*����4��xS�X�d[����Y=�^�g	M���?Mk�8S��Mr�o	��0�Bo��A�m֍dw��3����1Z>3�w���HLb&g.�1É��>` ���m�y�wE!2C��hklm�f`})�`��FC���ܩ��t���E��h��7OH�3��7��^���iu��ϟ��{XI�Ul�W'Ǫ@C�Cb+B���10TS���u����'6&b�oE��R0�F�Xk߉�y��:ϼ/Y�(ɋ�m���7�O�h��ګ��^L��U�x���,��ޛ�F�x�\ugЍpP�K�Dl>*��Z��=s��\��w�g0�$Սiox�1�`���­�7�L�"k�t5������%��B~��X���Ȯ�
�v�@��h"U҇����E����Zq�즐��ԲS�{ޑr��=�0}|��L	�`ȓj���[�G�%�,n�?JC�4cǾ��K�ߏ�u�,!���#a��sV��ټ-�<���=���6I�T����?ɔ�Tѥ�	�]��&}�j9F�Դ~a��Z0?i@L���&խ�B�A���/�t��Ȁmvsʦ]�u��Y��s�̚�t@���Iu������*j�#d�WRY�;�1µFW9􁞁�L|���Y���sz^4�!�躦��Ej�$�M����|��=� ��@F�Y�Y�����:�r�_�M�C�pģ5W�
�PjO�J�t�œ9\x�y� @)��W-���lӓ����^@�Ţ��d$��b[�ELpc��Ӳ�KF�b��eh�p��'D	9G�f�.�C	w��y�ų��N��k�L*����t�� ���_��`����ۘO���F�܉0��r���17ea��Ƈ՞�j��@<#�9ɉ:���9�^�x.���:#&�������?��o�7(z�A��H=��0�.`<)�����6������/�^��,�5��DXy
����n+��mi���{~�bB���h�H��X1��@	��<	�[���Z�>���Z�d�(������t$�f7�ՠ�M�A�.B�g�Ӂ!D������,-Y�!��Im��	8Yx�,2�`1�9�e��﯐����r���ݷ�}� ?S9	�(k��U�;N�C5ϐ����Č��EX�f�
9b�%���d3��R��M���S,��*��78!R���g��<��r�N�n�h@����w�#ܩ{x����~����� bK!���w��v��H!�VOm0�m����]̤I�2:��[~N���2������|���J��I(5�Z��[�'B����?�̱��A�R��`~�,Ú�o���g���HM�wn���`ʪ����:q�@�&K��)T��0y'�W���O��[���(M��>��uM��5�`�DV�P�Ox��Y�ܬ��Q�����;� �"��<~nQ؏k
��mR�����$�iA���K��y���Y[^4��[�D���Y�?�nJ0�'���	=�Q��,�;5�)^�Z��g�`&�Xz\�z�3���iv�σ�K�N|W�n���b��
_>r	�<n��t����of�a�h��x�Gy�O�$�E-D�]�4����a�)U��`�՘i�/5��C�ͫ)2w��=q��X+�rA"�Y��Mi�U5���/f�P��(m�^r3��q�u� ��cظaU-�$�|��*JZ�ebÀe�Q�y�$E��	�������FFa�~���_@��礠
r�?�HW�wΒU|k���L�Fc��O�����{�:!E����X� &�ߜR�'Xu�P����|��q5��otȘFVI�qrmܿ�Bc	f3l$����"�����W��?�߬��"'��0,���:�-�Cr�	HBK�3V�}�Ty�{쳁\�^�i�2�������֌]���o�-�~R�k��k �V<��������빚�I��}KjZJ�=����L�>0B�U��ɯi)�=���u�����#�%�Q0�@�)��?�
�p�ݎK/c;!%l��"zT��M�E3�*�r8WHΣ�+|&N�owUc�/�<��^i@�˝�Z���T� ξw��o�J��+J�ab����ʼG("���[� �F@�����B��V�L��Sې�	�ﷳ����2������O�9�T�S@�h*u)��{���φ(��1�a�I�,J����{!�=�yJ��EN�"�e�W�R�8l_���g�݅��&5HY��<���=�*�U�m`��_5)�!1 �"%��r��.��{|\,E��9õ�-繝��3L_��Z��E �36ݦv�y͝��2iCH�Xށ�8�c�I���z��S���<k�$��"��ƕ���Ϲ�B5QIѭz���R��ay�l�x/M���6_�q�^�}nm���F�q�C���2-��dMv��h�J�_��[g�@4D����楮@ܜ�`J�E��ա&����٘D�5� r �I���ⰹ�yFđ�:^Q:������}2�{�V��f :��}Is���8����r�)/.����5n�Ni��|���	<`}u�6R�[@���T��L�<���4�M��L}ܑ�!�l�/k*Г�D���[O�uaV�]V$G%�U�d7+gO	]��!"#��$𵨶m ,�*0�I�Lq�"!��WW;=F��p�b�BJ�%͂ �~j9���l�c���q!N�~ol���N+�X�
ٰ�S��
:eқ��1:"_�$Uϰ��Hx�G�W`K�cC���]�׎B�x��w�#ۓzbༀk����n������墸��\t��%y�c��3{ō�5|x�T�j�|���^,�j?�X��Ρ�5r��C2��j4Q���u��s.��]^(à���ܓQ�����.�1�˷й"��$�N�gW�8�p��N0�y�g�%�Zn�eۡ��U���Ӥ���;#�����~����`��S�v���qoQ�	��K�3ר��y��>\���Hf��P��i�;�I��RR��n%�Q�f�Ou���l�6�]�)�P�����Q˔� 5]D>��;�M��~Cv���t�]�zh���{q�����/Bpx�w.Z�_S��GL�p�Ո>�m	q@���WEaL���(�i��
6�/��^�R26�_�UA4˙`v_""���qF>{]�zy9&by�]�;����PqDȓ�9����AWЗ%'�o�q�f���O�$^|	z_�p}���u�J�5��{!<Ǫ]�z*���R㵽z���Q*|FZ�����b�9or!^P��f`������O��\���E�W���=�N�ґɨs��r���ޭMs.���7A��.k�#>�|��O"�<)Yx������T�
t\i�,bbB�����JX��N���0w���~�cH��g�{5�n݁���^WM�u��B�� �����QZ�R4����_���@�Ik�_�3�%��ϟ_������V߰!^�~�62n�ƥ��#���Q'Un�-�'��m�#O��`��܋\,[" >X��/j�d?���A��g�^�]zi!�����߷c3z2��'�"Ev�MO�3��2�|y f�ͳ��Co!��Μ���k��}`y��S����W4.F����<c`z�Ћ��j�X��,̞��Q���
&��Rݴ��g>�'dO���(�\�F��婹�x?I�y�2�ܥ{�T�F�hv�i�j���oN��ݹ��;����ˆ�#J`Ј�^C���-\VK��h�f���-�kr�D*�#���Pq=��M6ng�nʸ����?�.N��T�/�N4�j3�$�G�N��ibr')��Vj�s��k�F�x�.�Hog���WdX��l�D�֍����f*�q�>H�x�6�� ��M���O����M����{mU��#6��d��!��\���{��Z���}�X��G�jq�"x�y���odFu+���f�9Jb��C�0�J
��h�iʬ��S��?Ϧ���u�^�Φ�_�w��@H���B	ڝ�m�)n<-���_h<s���f�\��z�7ւ��+���7�o�s�D�m'@�|��)��@���*0z�C�XK�دWe����</3����
�����+9�E�/�
h���ԅy��(�r+���6��&M�d}D|3�$,��S�B%�������A����
�J(tbcҼ�+,Wf�H?.-rg���<�M���73���W	ѹ�����MWm���6z�+� �ւF
{h��7'��k�<Q�"iz��sc)=��wH#+.���jQ���X'N_�S6M?��sPI?�O�����r��҈0���ݗr���~�TR�G>4���/�)���cɫ��,N*׺�k�z^��msp������ۛeJ8p���^�"�I� ��VE�����AәXW���୔��i=>Tǐ[b2��$ln�b��Gǖ<V��_r�LA�2�؀^H�J]T�׆����y��NQb�:�������%*%���~6d?�ͼW�����|j?Oo[CV,� i��I�B��6�v�����\�iI5�}Ϥ�����F��WZ��Z�!��G�������P��H3��$���r�����Ȟ���Y%��_��<�@��]��^�����f�{��x�,���}��LADQy��74�	c��ر���e�!`���t�pHg(	�|�<��I��]{{��l�F�wM��1��ю7�(���A�m>�A��SO�a,M�N-�	X��7�I�xc%ŷ%�q$	�Y���PX
`����)X_������DǞ3'�P��u��R�9r�dd�(8R�?'N�!g��Y,��eV�G�ܬEJ��2&������dp{WsNa�B��EJ-,��3Nmo�;�RY�D22]�=U���tꪬA��H����� q����X[Oz}�nw	�	�_Q�U�r
���3 	�%h��A�g��Y+dϩ{�����n�s�����v��� �$����g�%'�EmJ^}�=�nث-����4�7nz�r!��û����x�c���V��5����Q[���2���l`(t	���PFמ����pBi �"�,z��˃��["�K��'�762z��A�|�bv�@����z�U�����+y��?b�ݢ�1%����($͆��<>���y�<E�� d�8�2^N�2T4�1�\A�����%��H�B5T�_S���}h�`�M��lӋ�aa���)��Eԡ^Hg�b%\w(��(���(	�ߘ����ӂ�|Jڨh���s��m����p`1�q�L�v@�D�m1c"@��Hn:^��G@Ԫ\8D�E�H�˾��YP4������J�9��{K��N�PO��������2�a=x:�T1	��k�*�����|�֮���gǮQx��xH;rF�l6N��Mt�:8�0L~e��1BAQ=���צ7^�)E�w}��><�!T@齑�띧�ӟt��<l��%�M�JF��BAs�ʦ�U��Z��<r�{��C������c�.�hq[VrV�G��t\Y�t��U7��fq�h�W1$���x�pб_}�h�t�����q��<��Qn�C®��?�5s,R��u�НT�Íl�G"�C	7p�b/;1�C��e��UJ�Iؓ
,kəv�1=�x��w�3.9��
�Y�_AJ��-���s��b�f�4���/��/P�7АL*�����vx*w 6v���w��!?1��9A�F��������/��U!�����V�ux��'��*S.w�3J��y/NSS^�����_q��ZǄ��֨o�k��������M�l���j�g���}?��/�]U'�PC�~��^�+�o\s�R����j�ߺx$�{�!X:�1����E����}�LiA���ފS�Q��M.�&`ND���n`�4yڂ�:������6��D�Y���wxR��Ÿ�Է�H�F�軺I�^�׀��t�GJs��v�t4vOR�������e_��4%�a�r4isĮ�h����y�3�g��	s����$��7h�r?���k�7̵�d��s
c�����= hB���U�
wf^�J3�U(m}�e�Wj�mm���.+wy!Z�4���|̈́�z�5�k�zp�m:fK�u%��س����%dg�P�#�	ֹ.x4��\?(7l��e[���:a�
�kѼ����a;��E\R���F{��Aʄ�7o�v5&�uͶs|l�]�	(�rAn�~�R�F�r��Cf�[a�}�)g~�2�w��H��%�4��K��)o��;��m��&ߕA-܅��`u�CDZ �IU�J͜L�	j�R�hE�� -���18u �E���ՠ�[ )m�����Dƃ9v	z��rT�"Rq�̕�����V��5 \oh�Q��Vl���N��A�f����x%�`���f�=�+�I���}�T��m0�os��ޜFߡ����J��yμ$�=j����!
��:��JZ�0>��`}W	%c4U%&8��z�&O�� �$<���߀�c�46j�g~��[�3?
�������21Ȕn/��3�
��FC���,��k�_7���� '	U��� BI�4͊�T�S���������7B��$�h����>�T䌛ThzPב��:�z� ^c>,�*��e������,��FƤ�td�^�G��9Ơ��)�@˩���g���>Z��U���u�03q�3��q_�&���>l�����	��Yu@
����I�Jĺq
��L������:����y0	9{M&Ux�@8�	:��p�-֠���lf�-� �!���p�;u&��s�'v�0�l{���lrOw�@Y��h�Ao�5�~KnrǓ*+b S:u�20/�Y��p��2=��q��L�?��{ܾY�?F{�j>"#��-�nu��K[�Y���/�d� ����s7I��T��:��&Y�q3�r_#vbP�J�j�]���&-X���� �H�M&H�\�<m��-���� ���$#�q�p�E���	R�Q&��8<�`D�s��f7l��]C��u���kG�aٕJ��Vf����u�?/����4gr��B�iU��=��]�;r�u=a|	֙�II>�Q�I���[�V��t`��@o��� z)�L��DO�V����١\lϦ���倗���Ui�����r.R�#\(�z�4�8�%}Ѥ$�K&�F���B�XK���я��v0� �R�`�Gs�3h8�������ߵ���*Eb}��������F:�+��{'\���q^?����\۳:��T�T�]W�Aq�,�� G����9ޠmxɦV�(�I���]�)�����Z�6<�����U!��1��/��
W�d5t�ha�-�>�^'a2�xL*��z��+YE�@N�Y[��s�|_��A�A>�{�b���>A���o�"����wN@`;h�<�e���}�u��]�7�/)�m�,a[Ǽ>���ٿn�ԍ�c���d* �5���TW~#p�Iݦ-���ۯO5�LN}�����"Fb��;އ�WRL���X�x��k��a��l�J���н�ip�ڳ )s�H�.6��ܟDv�u��kOi��}�e%m��q��~�D��3�[��w��Q�Ҋ���]��!�������4�4���������B�Y���̭�����~��#9vr�L :���r�@�
��j���%��9���S�����.Δd�(R^\��	�����XMKk:97�
��x�V��Ŧ����I'�YX]7�;�9x��^/ʒ�d ��nJ�5I������!r�K� (��w`���bi4ȑ��me���;�	h/W�;�xUӁ�����6�Q�q�d�Ǵ�m���b鴦�WYtgkI�2�Ҿ�7袜�Y,�xt���	 ���FU=�N`����n�Uexn4�xw�(�͆��M\\���Q^UTMt��
���غ����6{�R����}v��)E��,V�g'�
��g�������եr�7"%J�,E�.@9D�g�b����v.j�u5n��4h$m2գm�:_Z�X y�E�����(j�9�X�&i>u�h�M}�>�WѪ����"A#���4�L;��f�I(<�u~7�A�a��������c���L�%bT	�c��)4�"��=_��EMG�[��V��M���X�#\�J��>X�0���j^����|�)mP.0�@Lړ��8� y�m}݁�cx�=��뺉s�І�	dn����G��X9 �m�����AxsW�N�y ��WȀ5B=
ʸ���y��Ҕ�XR�觟߻b/K����:��ytf�T&N�T�B�þ��VD)H7���?8w�9��TF���h�<҂�žaN���V'�񁒠�jǐ���1��
ʮ�-^�nB��<�ԫ̼{�-X]+6H�=��Q}�G�}��*�d��Xd8�ªzk��b(E��`@M����f`��2�2F����I�%:wd�틍����(&+���#�SZ�U(����Y����������{�h.���9��;A Ȭ��Br��q�K� �r���ģ+l%�d�������A%�V�_��B|��������ŰYG��(�P2�߄A�E3�vE�k 	�-����O�� qʗ�9.,�wjMc�� ��8ln����� �Zhv�6jnS�5�}��r#ҧÔY�P��K|*ɵ3��U���fqAI���N��8�GY�� �
���#�m]5+�X�0�M��TxO$4<8�ג*��4zI��6����N$b��{��L`E�m�.������c>��  #Ws��{���q~(���S���]?+�va*&��v����Qcd�g��m#C;k��b��2�����=�Y����|c����x�yJ�G���9F&C"���1�Rן#�H^��ע�<w
�	��TD��
fz23����Ӷ]+����iL��|�QW(]�S`_���x���?#��c<��s3"L�
���9�W.�c���)�EUTr(u�4�X�-iF;����e�*8�����2��F�\�ށl'�D��*UQ0�'�$
���˚ް��t|G�	��c'F��P�Ͼ����݋/�-\�XO��J�#��:� ��5�쀳�&?bh�{�7�w�t�>����A0V�ݼ�JA�S����}�8��Ԏw=��J��h��ڳ�K6��[���ĳ�K(��oo���s��
�;
rm���x�԰������_��T��ٱ���Wq�T9I=�n�5S�Q\��~��K�x>��F���X�7�eG��ϩ���%ؽ*�b�l�@�8=Ea��1�6n�hOE��ST��++�$��vrO�����5
�e�d�#�OY�0*ms��CΦxy@܃/���צIQJ�T�N���Jl�F�����
vm��Kۇ�>I�>E�v"��c��^��
��E��&ǧ�xF�~��@n%���姰�֩�0����S�λ���~��JZ =�{(��W,��w,6��W��Dl�"ÏS�����ޱ�fU����mĮd��'�^fc�%����&��P�����.�7f\�բz��4}�ʅT��%�F"�dp,�p�6%��-Kd�U���M-�O��[�̍�!G� ���~X�w�ڲ7�/�/-�?�/��n ��.�sC�ߒ���C,6g���p}Dt}�(t��}�,��^�"f!�X�s<;Xg������<��8�gS��`�R��~N�Zv�豄=�M��/�k�M���G��`�c���5�f�x� #GuU��xc�d0E�&41���[�?�ւF��������㮯��ǲ�U	\���ܼ �fp����z�W@����q�?,�Y���*74�n���ɼ>�v"ܠ�uG�����D��v�2I�t:�KP<-��z�kaI[U  A��z�G=�w�25��K������L`r����w�	\��7|��%S�����|κz�2���7���Z�5���E��1b;4�A�"U�ĆwB� /u�t?�{�,����oWv=��T=��B�%�8_��&Z�au��[u���7�(�'��l'E7ݘ�:Ė�9to�Ҕ�DO���툃>(�Z�$:���ٍ�bu۞iT}�I��z���yt�����b����cswF�`X�()*E��BU�GC���q�M�rn/DFB�k��i�R�$��K� �@�!|`�z�e[�L�� m$Y��V�n���q4�x�_�p��pz��3��/��@����Eʫ�ٓf}hι��O9��.[�ъ�h��,��q�����v��z���פK�~�%3{B�vq����e0�iJ1��Oph��jؠ�.�.	#A�?Q|�I��lR� ̹m��^SOC�<����pDat�g��ضTmt?��o������
�g���i["�Y�-����$�a�D�X����O!��S�&��S�)���c�b���\	ư�k�=��^�GqX�V����Ӗm��-D�����:�L_X�A���d�SG�v��Vvl�B��$IBh��t�]��@o:��-�gr<�r�!H��:�&�<�T���¸dʠ���m�?��O�L
������ls����(��)�p��zv��'ZK�(�%�,�)M
�W�1����ȟ��Y��n��1X�~�,P�����O,���x*^�D��_��8h���/�P薀�h!-Y��w���v�߈Z	�%���!�]�]�� �n_`�TQ��a�N��'���MU�/8=B�Q�5�Pn������@��qY�_ץ�t����臑LQ1��_�s�3��V�����M�NU5�ay�m��M����GJ�r�8�-�Ԩ�9�r�/�б�e��P�J�Uî�i2)����{F|	>_��홉��y� �im_�ׇp��15k����:�i#����\Y5��h�nn�$�&�V7���l:h�3I;!:�C��幂J�T���QpVV���o��:�YZf�S��c1<1ї�����R�7��>\�/�������eb
,�^]��8�J�fF�/��j�vL�D���im�bW�����p�8%"�xE���ۜ��U�9���&TE}	$|�=u@J�\�+��;�0��ty�Ez�������V&z����6Q&�d:� -?�	2�V��N�p�`h��\���o_�6�eA�s�H7fG��1uH��BAP�a�/P��Д2w�F��ۻ��������&v�w����ձi?.)��4���w��ԭ7�q?H���i%W�׵�A,I��Cr��*+s��1�O���`8LʏV}57��ct58Ӆ����#�^�-Z�5{�:�;LU66��tvzo�8����7j=Јq񾇃�z��$�̺u
�c"����mP�5��X�O�gw����������WR�L�Fw��%���/[/�	�6	<��~�#����"f8�6� �%�C��K�ez��Ag��gfI�*��5���\R\ߛ���Ӵ��u�J��`����sƱ�J٦�����]-v�@`� v��W늋�Bl�a8�0�r�a�-,�[@ �oo��|�R���)S�D�x�1��+���FLm��&�q���a�l.E��-������]�j��$�n��
���(�p��[�d��N���c*AԌл�D)wR]{��Mm�j�]jF��v$>���+�y��K�;��4�Զ���c򛧬�@?�gƳtl6��Yߔ=��7�>�1P�A�4,1�0����ۭ5�B�N�����VddT�'Q��l�������H'�\=�nH�� �G������r���m��o�P疲��mD���O����Ē%����^����\b�����-8�ς���x(����8iO�<��:%.�%z�/��KX�F��k�R��*��F���-���i�s�Tîo�0LT���Ȍ@�>!�]�ў���7��ۂv�lB�j�k�^��'}���Y�l��������f/�R>mG�1�z����j9�RS裛����Bk��b�N�Rz�o�o�����7jm0]�]k�C�b��{��t�� ��D���������:V��{��L���E�eU�����L_����(�C�/KN`�}���)GS�野 r�͞��ћȨM�z��H�B�ܣ*F]BOyS�%e:#Kٲ�H�JLSEc�L-�3���
�OsZ�N�9d�m���q�5�v�������Ԉ�sK_lP�g�����,�/�!ԃ0���V��Ҵ�����P�+	^ٽ�i�z�D�	��^���g��ry~y���6K5ӣx�����H+ԃ�C状D�&6IK�Sڪg}�sE�>��Q=v���l5m�;�)w!ұ�ݨ�Q{3�6��_����D������Э���j��]�n�Ҟ�� Z���lb����.�ȕ{d�&3��B�ƭ�w�c��`y��u�z��,��sReqD9���W�v�k����yAi*#�"��)���/���:s:���'���R<����j��{%��ϊ�������
�N�^$�KnɁ��Uߴ)!��zy\�����V�x˟k��1:T�i�g����ך'[����X�0���WD�q�����T%g�%C��Dݜ����jb�2N�{/��H��|��! H���E'Y�n�qw�	�{y����bұ����6�������ǡ�U�F+��L�V���.�P��<�q),����hD<�О/&L����|�3��L:���}S�}���[V`R/_��d��B�.�'�V{r@�6����	��ڶ���N`��������N�rp�1n�H�LF�{�rү�p���J�o��rP��J\Fy�Y4@
f�o喰v�� 0���Ri����Mr�X#%��4��e��3H�-Ro%���_�Nf5u�	8p	���%�{��#�"��f)z����&��^� R#�u�@��h�B��(F,�imE��,5��������(g�.�#�ق�dlk7��a�|����t�[A��R�Ll(��F`Ku_@8.z��aXRf���Uj`�ˌ��T�N�U�l��&9�TI���,�Z2�;9��݃��d�{T�^����!�Q�_k����
�ոSW���mn5���A�]NuzA$3&�-�˧8�u�N���ܳ�|���Z�W/hJ�G..5ϧ�L(O@1�EYfķT�LL�8ْ�Q���cT@ht-�%��z���y���t���TE�h�PDT��~���T�?�Y��n�[l.Q�4 ����&?��	VT��9;/lw�n(M�� T����i�p��c0n���>Y�68Yla�����%���sq=������>��_�N��r��5
I���H@�-e��E�$[lx�Ǯr䤔��aCg�T�G���	�������|�߱7����8�h�s: ,OO�0'�=�A��&��!Q�ꇆ������6���6hH"bS�H�Ů�����Q4��\�f9�
���7w�Z֐x���V��3o"��#���1AIuQ�����L5T��)�6N�!���	�J�J� eQ�ɯ��l���*U-|\Q����b�ǘ0�A��ؓ�,�Ɍ;c��ݝ��M�}�����ą�in�����$��t���������(&�f��~j򺞁D&@��-b��f��|l�X� ��&�����@
l+�AΒ�V{J�m���ӝx�{�Eҩ�F
���[�%B�:�+�q�m�%�����6�D$�9�x��E��KF��u���9�k��[�����b�N5���	a�vD9}��`$s�^���{�S��a0e�k���d''+q�f1�(��r���rv�&�^׵؅�����d׵��\C��QZ.�	
%a�QM�P���g��lfSK���E��YjX��_V��'�Վ���&�x�(l.�D�����'v���u�^��>��e�V�c�z/�ҜbB�٬T�p�Q��ȒFv��J�b�3XS0��x6��Et�V�kh�S}��e�4]}���Nk���uO��D;���F�Z7;Z�u<����-Ь�����ć�m��*�EP�o�H4��t��9�A�r��;ϛ�	��n=d=����d�ƱN�m3�zWel���
��ㄭ�'����F0�C�ĩ��%���wYI����E�jp����O�ƂiSyr�wh(���wy�qI���D����De��0���W�����.����F��c�2�%�ia�_Ir�$!5�0�7;��e��s��Ғ|3?� $�W���1T_l�!Ϋ�����{~ک�Y��f����ǝR۩� �����\66��9�`��$ؽ|��{(!2\~8@)uXã�������.d�b��1�:�P���w��~��/e�9���n�<'��;�*�Wg
A�����H+ ������0��	���f�F�h*y�r(�r��Q�4p��Y�7�f�њ"�!�S���0�@Q`=���R.-��vs(�R�n��=~9�^:��V��^��^���h�Pvn:/���tN���&=�,+Z���+�;N��mG��2(�j�n�S{��X2��^������0m%l+�R73}`簰<�R�W�:��y���+��@T$�р5�m%'*wc^�;���R�Ƿ��D��-nhU~�:�Ũ����NwwfZD�|�C�~�,*�v!�^�Hptuu+t�N�VX:_�AB��D��
�d����Jm�^MŁ���.�w��!2����<d�1���t�9��:�L���2~Au7���ϛƋ�YO��!��L����$䢽^���G���M$�
2�� ?h<�_��iq��z�����Jwg�^X_*E������+aP`�븅�A�w$n*��P��u�ɝG@�=�� ~w|勢U&�ʈ����Dљ�V�����O~��^~��M�>dK��LE���\��h�&s�VZҹ�	�t��,[����\_�ua��9�<%T��Ǵ��i�E%��+�o-�m�Z�x��O;��T`>���2�گ&���-��=�s���҆���:2Z�eE��U�q�@]�����gNo���EO����'�����)2ۺ$>(x��l�H�)	�$��31g���Yl=����a��|��ؿ�h���3����������^)�����5�Df$u��o�|`��Ca�0���.�l��,Z�1��+:���L����3�=�b�����y�0����H@��Y%��l���������HNB�&~γÚ��ѹo����k\���x6TGTB��:9G�����q�!t�;�C��s�gkQ Ѝ|a��P��wd�QS�v�e:�ϔFѬ��^A*�]²_Q���M����nd�Af#�_'�Py$��	yV��M����B����_q-O��@hq.yy�Hxb�@s�X���Q5̣
��� ܸ/�:Q��g~k��2�:��qT�h�I
�8R�&� 	�e~�}�{��0݋������ɖ9�&��p@�$<���_|����m������+,#��}����8�����섫�]B:���y���d0��y� ��:�1rp+#âG ���T+g!7��ъ����K�L�L��g�Z�Q$���BkPs$�U-���,�\Y�V\�[Ĝ4!s_��;��%��_�_�m�3�-��h �?�)�JЇ-�i�=��Ei�O�\���u(�|�`�n��٩���%p\�Ր������D�����;wEU@h�l7R�Pr����e���w���o k?pn�M����0��QLO��Kn9l����i�h�M�J8d�n�C�s(3��)k�4et�8j�Md�:��W	'��0US��K ��e������ߡ��S������,�+���yaK�R:C�~��SV��m�2�y��1�O5���z�<% i(��MԦP\��˱�B�g.��7W/�e��s��-�[�:�<c@q�:@C\t�|�W+Ƣ��ԯ��2�2�y��{d�[����D�FR6�"�_�.�����D')j�sk!�� �>K��_6���rظ?�M��|0V=*�^J��/����b���|�૽�#P6��	Ǹ���c���IQF�D�OƐ��ױr�L;6�&�V��n�R��sU,��#�!�^	�ݲx�*�z���m����D�
��O6��ױg"AZQ�>�)��*a\��=��H�ʩ7�ǘ2����J�;רM��0����cKR.�%-�R_�|�Ƃ��,�IYS�SD>���DJ��T��EieX9F�KV6��M��6&2ᰳ��ґ�9w������� }�R�Ĉh����<v��o>�xB0�qȆ�����,B�`����'6Ǉ��8w}Kg�F�Uq���:5?Vxu�V����9P���h�B�0�{��L�@f��
��v�� ���a�Eb����,��b�S�*����@����b���'�Hkږ��)i�~#���si����V!�� #�����/3/�_��<��E7c���!�_uwc���9�	k�rE�	��6$����Q6�a�X� �a|�i�ܔ�I�h��	�}�FD�u��7Ʒ��g	A'�Œ��;����#��ı����	f��y�aGs���7QK�~G����֠�r���+�����>e�R�J�1�nO��C|㼰���B�T|ޖ��^Pu+_N)r��RW���_1P��HGUf�x���?cw�8q
�	������BD��7�v#������*�\J����L�C���ٿ�.�r��=�Y�s>��l�*���A��rH�Ҁ���C7]�!es)$����+t�}i~dE�D�E�� ��"��2=7-��x�����KZ#�a��LEJ	E)�
�4�~��P?��]@��D�:�b��	)�a�=9��_(�n@v��q�-)��L�7����UY$@���>�-So/�?���SɾFb�xN凼�?�<�c�7�5��- ���M�_��`�a)R��WlA�ҿ�o�gb�b� S������௠Lj}7)�zcWq1s��`]Fk
��&̾E6�pF6�� ��B|�E=��Jbu"�υ��$�"���^L�ޔ��1��!��v[�k�.�e�PM�,�bk�_'?�e�1@��X����b7+�M-d��:A O�㩥�]xw�_|���\�t����݃M�Cۖ�����%���G�ueZ�m��1d�bɓp���)���^��u`��Q�(���p
�B0.��e/~�(��g�{�{���z\I��'�?o�jhRNo£A�G�N�/N�����31�&��4
 �Y���_���l��V�2+(��Ĺ�"晇̼�O����*�Z�j-��X��Л�/����%�CI��;��`�y�k��G	\����N���ǆ�I��j���\#�j(Ȣ;�����%T.�	���qt��+ �D�BOc
J�,>��
ts�{���\$
\i�q�DT��ޤ�	�:��/="ᵉ������9go�	h��<e7�4���iZ�px�o�/e��2��qZ�eb���*�~���U�Q�8��9�Ӡ��>n^��{;s2|/·P{I��NֲU;	6OU�����&��fa$6]ڙ�M!k�� U�[��lK�<88V�J{ n1�Ј�h�E��<�ʷ�͎�K�Į�"2{@��.K�y�c�%۠��e��(�q�1B���&3��J"K[�d�>�@0�u��º���p|��匓� �����K��|u�vB6��鰁!=uY�R���-ں�)s_G��(�^��Z��a�`頖Y���[�,P�DƯW�V!�oE`!��Py<97F�v�;Z�~���`�2�Q����������m�)�iC&{6If$���#�6��͑�Ο��;V~��NR�g���W�Z5̵���H+v���a=�B ����cߣT����>�+�W�x��}�[/��Y�p5���{2��	f����c��ɟ5��쇩9`깳]xf	.�h$b �a�=	����4�޿���7�OF�f,o�S-��m��_�h�Jit?Y�\�h����*�W�ukN�N!�b����Y�1��>!��f�A�1����)�kk��%6;��1KYý�@}QM�9�{�M�Ӕ#���`��4����Dw���`+����(�A:� {eǱ{|3� d�=��c�NBj�'O��g�	9(��:5P�$�=2B�y������CY`��s�n���CPpVv��R"�����<FUn0��(b�����!<�]m�iX�tFܟ��x^�Iq,�+�"6ށh+y���/L<�Hq��M������_����1G��"��<��� ����@�5j�w�7����!�`3�'.f?�Ʌ��YOJ�[a&��]r�J6�2+}��o�lL���x�$��.Q{��Z��U���w��\-,Ҡ�v<�S�1�]r��TE�-��جv��I]��z߭nA���{Ӈ�l��߹�Ͳ��V���KvU.˒:(�NiW���	���B�d��>�6��|\�k4�"�`�Ć��5�@7��	�v���$���t ���x�vGiӣj�^�S���[s��FN �q���y��:�T�c9��
\xG=|$��i�`|1L�L����[��M�2}�"���G<O�vݍ'��E�����C�+�Y�'�plM��2�rB�z��hU����F���?�ԩ=�b�-���֌wH�H9{֒��?��k�~�5��ߓ~|��#�i%Ǧe~:K����"ȕ�8	�����P,�����)�͑ND^�}<�&&�c��f��Or#ab�O�5{�Il�Y���~��046\�����GQc	*J��NN�Ij���.����RM�Ùد8��5��6���O�E8(E�a�B���3$4=s���nRM��r��ys����B�ˎ�zI��]����Q0����:����A
"[�9�������n�����>�Gs@�E:>��:z����3D����HO��F[�UZ���L���5�{öb��� �Q��h?��d�W1+f����a����]ڕz�Ѽ�(�*�
!'�^o4v��j�w�s��+�J�5�x_rY���6�Y)��PN�Fۿ��fΒ^���;�uJ�+��V�І�\��I�~/�x�,�o]�T��{��W��CDPw
7����K�V$�U�@p�O�I��V���eĊ����dx�hAt�q��&h>K@%7&��'J/EH?�ȺWI���ǰI��.�V�	�-�&=���0C\��t;�	^s��ӛb��F���3�`s����J��QuG��;0�ե��H@�{�����W�x��|���ƻ{޲E�^�%�#K߮q� r���c�d� zS`PKi��x���`Э-�m��(5\8��NI��̹%���c<h����@S��d����־>�F��֌��=T�;^1<�4#��x�a�t�E���I��Z���͛����*�!3�	+KG�p��3(����	A0%3F=4$��/tS'xi�L=��vBP�z$�l�7��7l �at��>�;ީJ#�����i����I�rٵL�ir� ���]����u-��:��=�P~���*0��⽴��.8M#�
f6ٻ�;魚�	ٵb���F#�:=W���45.Ml�%X���tZ�؆-�������oba���*&`�D�Ĭ���(������=����;��"u~]I [r	w[�)��0P��f&��7�]�]���UPs)F�1з�FZ�����
2�_��?j���╿�`l2̓3|��t�M��s;Z�;ot�x����V��(I�� e�s�PĘ���üH�?������s�sU��1��pҾ��oܻmR%�i���Nx���o�1H�5.��v�e�� 4[?��L��F1�䃧0�!'��z1� o���nݾuv��-g�y,ٽo'�0���M�nJ���W<��H��cH�`�ti�ʿydM���3SAZR�ѐ#��Α����zI�����ve�'�ɢxW�����0�c�A��Z�B�C��p�����%��)���x�\�L3/sd����V�;��~N$�8�Q�A6���g�kr:I/��OP�\���b��U,�Jw���q����
��T�&E��������v�p(�k��P��H���'j����jW�\]�B�� ҽ[z��\ܼ9����"��"����L�+쬕/G_}�>���QM���~����&m���JP�ms�G�A`pjL�Y�Kx����  '=�Oń�����Ў� x��I�RH��e��H҉JDkj'5�V|�{�����XJ�#��~���Q?��K|Ǟ�0���3T�Qu'�hBe�t�֖�>�1�3j�3�l@���T23��%�-�C@��v�)�#����>q¥r��J�0?�,ɰ���:��"O�u������:����+z����A�.�+u����Ϲ�f�	�ܔ~�C��Br�A��f�����@��	T�O�\����� �O>h7�SE��e>���I�=~R������;�G��O�r�e�;�� z=nS���v�IL��7���{��*���^G�X-̆�3�ӗ2��l��F	�G#]���O�B�uYP�4<���d���%���:
a�!-��M����%����c�Kw��|+1�K�AG��E�c����d�2p�V��p�!��)|1Z���.��C�=����,�r�|���5@�Un X�Z��v �����j�ZH1lK|ARn�I����w�`0<��3�$��R�YJ���¯7�?4ʩN�K2��70�GF�N����ϝG���Z�W�_�������UM"ӡ��!�(*۴w�iQ<�1A��wǼ��<3��v%�D���T�4�y|X [��<�VY[�ii�?3EYd����#Ӈ��d��]D8��s��6^v���!S�X2ʽ�	a-�� w�3 D�s��j�;�O9gz
���Xv�٠}�7P��cLi��
I�'�����~��1����4m5��0Bz�s�>�����-���6������}x�^W���G�#Ѩuo�;�J��k���ZL�+[�3���]�+Hpy9�3����u����y�\"l���F��&V��Y�� &N۽�#���@�k�FP"��&�����U�)��>�ȒT���.�8��l	}ցӹ~Ys%�ұ".�7O|<WePˮ��}ZQR���u��C��v���ɟ��Cr�O���Z:%��9�8n�(��'<ˉwz���9���*�x���7��j;��9M�~��0(A����w��>�k�i�c&C݂|-0t+�>@P$pz,�qi�m'�R�!�SlM��p\�2�;���k�e�h�XR�PɄ�Xb���r7�!i�$oml���s�Yp:V�u�I�^"��v���"��SjLK%G�d3�Іtwh?�֎,�D[�t"��[C*<�Ϧڄs{��4H] ���]�=-�J��3(p@� ����J
�8/�k=��;�x2޳9Vi���xvO��f�y�ᢎ�hTa$L�uzLg]�
�o*$�==�#�.8�%C�%���-&f���R{���A9>c�\�p��[�c!.�N�����&�
:O�N�p��ݲ���2gjM�Ue�joH���!��x� 0�E�4x��	�i�LS����|���n�_�X�Ÿ0k4)+�
(�s�}�oV�Sʱ����n9aP/po�VJ�7�����i��Hu�م\0
�}qK^ �����<�V72q�Œ_�bv���*O��&+F�����E�#2�4u�mR�{��n���+Rݱ\��`Ƶj�/���]�(�A��Z<�7�Re�;�"V#�/���l���笻S����Ћ�����J���bA�3�W�Q�(b��s��;\�����	Ƨ0�"�.\�C����FW��Lm`�8;Y�9U��a��"ंT�q4�x��^�^��ꔅz6:c��;�)@;���>}��/�a�� g�6b~�,������p����@�Q$�A�/�Y�O��㑛�U6�0�'f�6)š ��"�x�`"����M<� w��>���O�x� z��ȮG$���k�\$^�>�V\K�Q��s�m`�'���IE���#��腼0"�u�����D׸��1z]�;�u:��,s����}����I�[�g�3Y-e����~�����W��١&���pf�9Ϫ"�MO�ִ�����3���^D����'I�L��^[��gRO��Ԡ����/@}���"��ƂF9�ji�u	���\�[R\
�X{�5S~YQ�gƥ���biu�9�|_ڄ�®��wo��1���-V���W�Uk��v�L{x�!7ET���ӗ�Ӑ@Y� uwz�0e29z 
�4��=&�T�8-�։ɼ�[�b#�0O�n���#$áR>�d�5�T�pn����/�Vye�&�}����䮀����KzD���gx3����)���ag&Y��Y6������P�7L��.�7a��S�Tn��S�9�Gk�����:X��|n� LV�].B��Ξ+qMC�������	L>�,6x<s�w���ƀ�
��N港��f�~�p�t��)����t�ܔG�+O�,��v~b1�r2]QnI���f��sM�`�N���8u��iw��0�ǰ�D J�2O�!z�e�j#��^�&�hp.�30^�[L�f�~���V�A����}���A(�Js���1畕i�RHX��������BT��o���j���栾O�=<��}W�wҾ,_:�pW�SJ�>�
aڔ������T��5D��%oֹ@�#]��'�h:�/w��R��vEU��yyi�ݼZ�,[�;���U���#P]	�moX�	@�z�����=�����,�~*ft*	��c�X�c�{&?�Un]���B��8T1c˻=� h�*��e:.n/2DR�;h֞��Nj~�e��9.H���i<Q�� �0܏�����:��$kO��q��9梏�C5�Ki�f���H�R7�Q=ƳcK�$3��dA��P6
y�db��Ua���zX�DŸ�UG������l��r���9���;w..�m�oe�vջ,�rbxv�J��V�؅��}�M���Z0�� �th8ѹ?�Cb��U3^�7I�ס�}�A�i����Ep-��(�#�)��v��k�.P]a����*����'�����T�eP٭�I�uY�G�ɹ?���yXMFa0��\�6�͉� Q����$���&[�kRk����7'�7��m�&󗑏a[Ԉ�u4�mx��W Ŗ�4�>��H�s޲��1I���ڳ�[ͩ��~	랽NP�?�� �{���;'2�m�'�M�Q=�.3aG3Z�E%[�XB��Ǝ����H�����PTu��`�[�(C���{��V�P�0j4���Kg�yeƬ�A)	�?�Rȯ�&��%�����W���A=��Z�����;�1�G� �V@�%(���<��L@��yL�^]�n��Vf9�K_7BA�M"*"e����o���ެ��h�D$��U0�f�Up2��2���AE��j8�yzP2�::j�!����[��|��;�u��Y�ɢ]z����Sʥ��0���y����I�PFx�;����q��"CY�B��7�V)�ko(�.�݇���(9�ٞ<u�[��R���sT׭��K`O�SX-i.���wO9��=)rOl���x_|�`�bw؜T�����p�l7j�%�\�����Dn��wFе�sO~"����S��y􃁬��\�g$AW��iV󿙸9����-H=)4q�*��-��`���i�.6u�4����;��\v��D�oy�U�m�p���A�92��.���#v	���βH���s�Z���O6��t5{Ve��vv�Go��E�;�(����Nm}:%�;�S�x�Ƿ/7���T���c!� O�N���b�;�L��Z'xgB���)����ʽb���N"M� ��x�䆻����]f��|0�w�}�u���K�⛣�8}��~2�G�#m��"�7ב�jŵs'�fp�q��?�t>8�l<P#S}���m�AӡE��q ~�D�����ʱ�f/f-��j,���W�S	����������m5Gtp_����P�)vY���[d7M�b�)��r!qtH��A��[��Gbu��܁d��{��$����>�.Uf\�h��Pa6��_6�'=�9T�VW]�^��E�j��6�F�$*�"�N�N��(�]0��@���虹�C���w�h%�Bp6Lhs���s�S�0������A���6RW��~9hf��H���~[2�Α.�װ*��u~B@w��r�A1�\�ʧ$��=�9�A+i���ē��,�Oue��� �}o/�I���e�8tߋ��)7ɈƤp�:�Vm��
�w2�w�x�ED�0*jg�GQvJx�(5^�:;�<����X��6H雞;w�m?�� ��O�,���S�� �X�=�B�lA��9�:�}(M�;��q�g&`H�e��謟#�Q�����g�=�B�,���˞R���a�9�h�M�ꆙ�ޞ�����i�j^��[�L���W�Ru}-t���J���!t怂k�����Y@���3�\-[6���8�2X�:E�ٜ^�I�:B��׈��|�ާ$qzx�����Z�"8}!����i�c��Z� '�XB�N��CM6��+��[%��R�[�n�b;ő���s�D{
6��	�~Qn��Z��Dܲ�|�Gr.k|8�x����>Gq�nM���E�� <W�N�M�ٜ�C�2�N�T�FZ�V<��Z���[�� ��'�b�.��r��U��8U��-/�%(�WB�oS�l�i(�7�cq�Ydd�Hv2��M@��%.�_���+�O��O\*�G`Mt1��Ŭ���������Ԁ��"�z��Gܢ�Evt<���v��Qd�^-�,�|[���ו�sۏ���>���^��#0��JR{�~���nu�/%:�Ʃ�S;�W4�A�#Z�к�++�#��*5<��P�I�z���g���w�byW�?���v�(.�G�.��¢M�"ˊ[���K.�9�Ģ9�Uj#OB��D�2��ܚA��\�K��M _<\P�z��2�uD;�1��ƅh�� O7x�3aw ���M��d�*,�K���s�i���9$���R���{��/�3#v�V_�ዘ�C���i�' E�Cz�ǀy�\�f�8��XFk��̕�Nd�%]}�;�S����<�I��./�Ot؆S���;fJ�^�����Z'`&�x� >�p"��Y��Ij�I��έ�$�e����H��UT�� ��:����y�r �ȯJ��M�u����s^P����s-���#e��X0X��ܘ�u�Ȍ˹��<|}bZ�0��5���Ʋt)�1Gw�6i�������S�utЀ�AP�_�HHo�x��� =�90N�u���O.?-���_
���+��E�&4h�#O�^����7`PeS�s���nW�Zb�|Q:{�iN�n�qs�m���d��}�̳oA�Q�q�"������r��Η��_N11�L�m�@`����:\Rϡ���F�Q�����`�q��*.��ݝ�%���4�&�n�4����l���/�ܢ�XV�Q��&�M��L��6��灒P,�<���*��ܔ��k�G�f@���~{k�}��	 �>9���<����Y����.�G�yp��{�g�@G�dj�v���ƽ�ю�]B�9���ibv����u��"�ڤcxj�-B˛�~)
�8	�!=�.;9Bci C�O�M6^�ڸT��u堕��s��LhDc��bz=��~B��s� .�7����XEJ06J�QxT:���`�0�!�)Ts���+�n�G�D��X���7d�"�L�j�B�"*u�N^p�p�h��W�G���&�'��si���pbж�P(�Ɋ��3�M6����Ƭd�os�hoEz�8��x̽ۼ(��(����Jm���4)���X_���/��:BVf 3 D��C�뷞X��$�£7�#��K��(7�i��]l��\zG&=��
դ�v��A�ț�C�C�º�=���q�ٺ\�ٍX/����ݜ�N��?Z�<�ԣ@	�~�l�7�����s,B���t��y�����Zc?�'��K����+�w`uΧ%�gB�XO�����j�ƕ�S��"�h�6�g�Z\��b�z�CLV���l�,bB�,5n��_Q�@2�Ym�w�3'w5h �
��:DCc�j���a���uu�
x�Fo�H���M��9��'�}B��	ʧ��
m�3Y�ck+B�F���R��ϧ���>�?��1+������}(�"��K�I�5A&�W�R�mq���dR>|�m9��Ķ�T��)������Ko5�r	#i�-$���oﲄ�/(����'?�Ll��Z�i���U�Hp[�!�^�6(�8gzX�oS�#����}E��Y�\�c"GKU���#�<��u����OE߆�:��9rL��|���"K�����9�����.f)�C����-�8�TP/n�Ȳ	z����Dj7���x�C� �1�1�c���.�΋�~�ð�E�]M�������]�XQR��E�X�ʔ�8-�^xj���Jǉ���ې���Ka�4]<�;~6�^`���@E�9|�y{3�Rk=�)���
)&BD��]��";=��&��¿5���a�S.dwC�����d��h� ��C���E�B�_vat���<����a&�t�r]��䧮6���=}�;\J�԰a�T ����ny��ª�n^��*Ы��LB\����_L��s[b`c��Oq�s{�|?�9%Zՠ��\*B�z_�4��1m�`��hu�K��DBf*68~�nl��dq+Ii�m	�=�1k�D�kҼ��i�����w��GT�[�v����H�(t�X���#%��E�h?�=�n��ғ���ג��/ʈJ%)Jd����V���q��$�2�t�CJ�|���M�:RA�5���z��D@VR��̹R(Yb&�7���M���e����z
�����]�7���s�����ZR3��{q~э1ϗm��l�skf�eT�͡@��,�@q�o�iP�g��c���H$[�'�ߚ0ӖPJ�������1��_��x]��N��$��(����"0,�,���e���ʩ����������t��:����j����A�D�3Y[�ȗ|}Q۱ #A��S#m�p��e|���ir<�m��x�%�Rޏ.�b���x(f0Z�x �r+[˰�j*��N�K�\�Nso֍�F��:��������4�-:�?�,9���֯F��@o�*ڛ�7�������D�ٯ��Mƒ��{6�$����w��m�ކ������os��(jTz�n��[x�;�i�IS��%�{�qշ��U\<f��۝ϕG����P���]*�-�}�)�i
č��?4ꊩۺM��]��e�&F����1�n�5K���=��Z�C��(��׼?�?_��zRi8��!�юW��B��ϻ5 h�21<v����F�;&��+����l�2
Ļ���Y�r7b0���x+�M�?L�ZSl��}(vz}�n�7�uS��M��6����'�wo_�Jښɭ̸�2�p��h{)�ŃWZ���A��k.��;�m�Ȯ��ϥ��6�tN�#�@���m��
�VX7�5CƉ^$,����wQ}$�Hx�`��s��+z��/��� �Η+{?��DŸf��/��YA��@�0I�&R06N�L��?���,p�)�%�R��fG)�f�׷�}�@�*)�q'3%��Kd�Wr��]ܟ	x�KW���ګ-�G���܎�2N!�M��3+	~�l�*�y� ^�Z�Z��!���c�;i�*N�ݍ��8\]�<���H��6}�2�Մ5 @i{\��ir��x+U^:@�|u��^zH�~ -UPX-Ģ6�c@<{�A��+��3J�����-6���
2Q��s��T�g �	!�?<W�0->�5����}H`g��T_J^�؟6C�A~ћ͛k1�����i��6#/M��#8��[���Ϥ���G	�����V�dRK�b��$�-5���[QrՃ%�.S�ޕ�e�8�Ջ	���VqL9Q8�� \4�d�F�!�&nL�U<�āK�X8�$�r$�_A�rir�E�xُ���h��1F�1ݜ��N���3֔�6��$7)@cR�V�,��\�c(CQ@��sYU�Է�1(�B^�����v���ZS{�M(���arzUn�Co ,���mO D �v��N:�;��b�����Ǳh���*BU�I�K	k��i�>+��A��N��A.���y�
<.6RW{'is���,9��~�b��J��7����wW$�ڴ�Y)�����6.����������s�I��m����R�Cm�fF�xcV�� A~a�*�:򱿉~����h�²��wJ�9���"�P��NB�Q�(��f��e��D����PqbU�jC?���*���K���6��y�v���=e�V����Ť�%�߀��ep��m��Y@l�f�ȥ�ʻ,� �k�7��NP��_+B�R���V#���S�r���0S\ c��S�����\���P����H��K����O��a�&T;b%`��~���F;xcyj`~B����,�4�w>�`�̻���у�
i60f*��������ֳ����~,��1��܄�o��	�|.)t��A�c0*v]*Vl|aVÍo��.�f���ͷ�����S��QWn���ޱ<e
���}{�x�hzDS,�� �K��} b�1p�É��(�,~�N\���p~���b\��#U^���?��ݎ	/ͷ�v�P��u�ۊ$���q :�C��[��Ө$�����A%�r�Љ���u���W�</�;#9��΢#��u�4�4]�n�AJ�8w-^�9Ϝğ���w\o�gT����L�P��`h~���/�7g�߭�t��K��-wAG���&�/gD��]�����5�s�i�Yer�UuW��l���c�;�f�%YuQ�
��%�4����:�y��e'E�]h��Ӡ_5ӓ6�Ep�vh�@�I��vr5��b>��W��.�?iO��������_{��L߿��JQ�2������nU�E}/�D#n��u�g����ȉe�Ϭ��|1��n�����e���QB�3O�|��9���H�z���f������j��QO	xT��)�G^���]�u��������9E��F��ϻ���3�V^��R3 |�mN��3�ܤz�=��#*E_�[ɔ�:�z�}���yJk*1f����1Y�;M�-|���H\��N5mT��y`���p���Y=Y���x��o�sٙ���Q��"��E#�"Y)$O�~"�O������~��#�ܦ��F.�����#18Mb����H%ˆBU��|����I���6�C��Q4���
�M���CZ��l��Ń�˽U�6�o]wp�`xU=vV���4�Z7E�s��q���"D��]��?gH�:▹����î�8�ȿ)�?Q�礥�W�}�.5	b`��ؤ���1�~l��Vp�:�K��_�_c�R���h�������4��;�q���`x��Hvo�4n�'7|a�����sr����|Sdl��A5��A�_�b�@h4��ژvMC����V8-�� �x�̔�����nl|��[�W����3�W��%�ٕ�x�8���jn�g?&�OSL�9c��a�=\�v2cª���V]�:j��@T���`�+u�Tx�.�Q��al�T?k�H,�Wxu5>��G7����|�~T��[�9x�Ebz����?�����`7��)�v�K�,�ӲS�o�4B� �E4�2��ť_plG��+b�)���_	�������������3���Pޔk0����vZ��b1-����,����ߙ��#Ip������םM<�Jd��Ҫ���	�oJ�,ɒH )�#7.�'��Xa�Z4���87I5���ڧӒK޸θ���"�%��"h�Wɿb���U��h� K���E��[�k�L�"��6O9|O�/�|�S0���5�n�?�؆-�=%�� �q��ߛnS�A����������[�:��Y��z᪠J8��n EꞶ��*��Q�'��I�|R��H8:�.�N��:��О�$Ǉ�C�v@\��Һ)�a#L�rm?�6�0*�9�bN_Ev*�B����k*����~��|��K�������H%�Z_��z_z4/Y"ۓn��6�M�#;R��E��m�C%ݴ����I_$��W~p��&��vl���9����Ǭ*�,a��.��-u&�T�K� ��	Ġ���5,�����5�~>s�w-I�C�k��'��>a�dy�K+�7&�l�M�Nu+;z�-[�ǁ�OX��h���+��4�4a����!�ܽO�6 ad��,��@a�د1^�(Ҿ��u��c�l�U>4U�5>6��ͧ�)���?�\Y} +C|��Fc���.:!���"̿r���B���x�qh<��\�{�:�|]8�a�ȁ�~�M�4�$Tg�\�tj���5��	g"4�#���Ȩ���w|��2�~���4���	s�F��G_��'���+�^&�1Z]�;"$��ږ�z�D��#��kI�N�܄�����>�" "��	�����}�"U�"]��ѥ?Ng6���v�lO�|�fڭ`ҏJ�^_���;������.�?W���0OG �>��~i�٦�a ������PN�c�t[��{Tȧ�}�w���#��k2;8E>񲻒@ǭPn�=?.&Nc�v�?
�3���"�ﰡ�<W�r7���K�nٖq�C��ہO��B��#�GUã4�pHR(�*b�A"fVM�-�w��&�/���� WU=��7�c�͡�����43	�KZ�>`�T��Z�)y9J={>~���ƾO������i����{�gUq~<�K��&4_E"��U���#��*�*��[���ʩX)In#�:��󛖳�'�G~�l�\o,�{'�=�	�V���b�ɣ�Vڡ��sU��n|~ z�B�?�b�^64w%���5Ui�� ���yڞ������F����yv8n�?|��b�!���;���|R�օ�Zx���F+�5¥���S�`�D���8�f�U]��2���=�p�Z�?N��-Q!�Q�u�m����t��i�AJK�_�g���Ks< �b��K��کK���M��q��<h�*j)��$2'�T�����T	����pEaJ�	�p���|+|2gxlK�kzb�z�\��k(��ߣ�s��?/и�D����̖pl����=�rxg�������ͼ��$�/�9BI��6)�r�}AA}B��$�5��gQ�+��x�xgN2=��bj�,�>���"HZ_����7yo����`Qn�Ȩe���V[�������۫��J� cdz����P�
рd��U�-8I��du�8
[J.2�LCN�o��Zq�]�w����g���M5��VR26�9�P��C-G+q3�w`}�@P�BO7zN�`~�6H\	�/r9�w�S��7A��G���y��+]2m��,C�	&�N����2Q�W�5Z0���k$8.I��pJ{&ߩ�N9�(�k�����Y�ύ�_ig���F�E�]�:o� 
�p�*d)�H��9�F��^����E�z=m
�.>z!g�p�ҽ�F��M�ܼqZ�5b�h;-���\��Y���>Ӵz�g ���jB���2�����Fya�1�2����
���*	���˓l3YS(L�̾_�\_l���e:�+ni�ʇk��"����E�ާ��m��n{��D=�Y�OV��`�Q"���������j��t��@�XL��yodq��ra^(���rdk�}�Q��A�"P��iVuej��g'PO�nL�z.�rR��&B�b�_E��>9�gZ�����$H�\���>DX����
�����}�
����_l�#�8 ���`�XY�wߖO���.Ey��x��7IP�]��|�v�p/��ã�<��5�n꞊MA�u�!x���/�$�T�qh
��t��tc)(_�|k�J����>8c`��:f?���+�q+��!X���(��X�����y��5��Rһ}M(�9T���f����8w�:_ad>���}����heioo}T��)��3:a���&�b�hy�%:МE�	�h;{�� �/"!}Qܣ�xeLf�*�q�1��9&4�/:Z��rQ���I��Э��P|j^���y\�`�}���q�8�A�$%^�p�d]��N`D�ΆX�䳤�0��N�m:�(��n5ezE)��k�8��	���5�ͫ�dF��A���U�
�V�y������W�3��?`�+���=<�蚨"�&N/�޼Y\}�ᬸp@ @�����x�$�q�w�)��W�l��;�Ri[zN�|�(Zl���&��*�pH�c�|Q�4}���@�Z� �7t�E���K��	�h��K�>�h��4m݀��d��l,;#z��\��%zu�m
��Us���S�mR����S�=\�X�D��.H��2I����AzC�}c�>g�p�B�|F_��g榡<�Gf����z�'��k
p�m�� �͆}�^'��i��.�0P�fѢb�`0����Yqv�xqyb�y�E	L<H���X;�P�q-^Q��#(x(�Ɨs��Èw�0�c�A�=��S ��!Qc�ȬN�w�)�+��<;��;3k�	�R#s����B�5V�-�uYČݸl �Jj����h�����\�A�����ߎ���t���3sʕ�¾�
�$�eu���mͨ����i{��g�Ih"�%eA��y�`|*�9ݷ,1������Pɱ��y��e;4�?�v�|�7��=@���k��ᚙVf$׃�3:����sê����ی�2)Ϟ���.(��ߋ&���VΈ���l�ȳE!�R5ǽ5&��;2 �7C���*v��(��ɟ�$9Y_Tk�:F(��a�@-�N�]zʴ~�����f���p���]���F�ί��o=�jc�d�D�J�����4q���w�}��>�Ôl.J�5��!U=&>���.w�p��nE��'�I���~�.��Z؁������1YqXu�t��ڄ��~yT���,0�Y�� �n#��{�3nl���D�*y��P�)��`){���?�SY� 4s<�7}�c9��[�]�������"r�9�NL�V;�"��r��4��L�\{�q��^V�#��[�ɯ�^J���˞�M����������h*.Z0"ؿxZ��­����}T��l.��%M�pRI>j��X7XM7^oA�7^N6�+m�%�ޠU'y�&�9������7)G��%����Co��\KqyP�KcW�k���;�~)铗LH}v�`�λ�y͞t���ś@�G[E�i�E,�Oo~Г��M���R6����~���S��oU���.S�m�'�9h
�J���Gy�8����Џ���w3��k��'_�H��	�V�:2
�׬���FĲrI����O��9!�	��ﵤ�'	o*�xJ/��2�)�3�['m��Q/���}?��=5;o  (��34X����-�@S��JԞѯ
�ڎ�C��:�>�2��Z�I��T�}t,B�>�?Ah0
@�n�7m����F�k�Yh����p?��?��L\�\+�W��*��B����&黊d�j7�d4�X�'��]�EV�9Jb������QR���`};Bm���7����ᥰvR�G�ȧ�j��J��\匯[��P�O}܊�c�a�ԭs,N��xQ7IT�b�9�v���9��9�V�Ꮽ�L��0=����!�n�ʼ�R�4ſEW���-d
�@��2�*��H��l�-�.-�DP�d9q��x:����[��W�4�����_��pC;/�X����%���DqY���AzE �g@���̲%Be�RT����l=�	`n����{<� �/����PL�[�����4����v<��詐�y<�0�*\��
�j-TI6o�^�A���	U����UDKt�x۪�0�@j(?�99���a4N4���<�TIɣ�7����	R0a��?U�~����������j�p������,8��w���
R9��L�)���~��'��M{Ʈ��֏s5���F���������z`z��kϾ��	���W1�?:XE�|�n�.M%��4�����;�����i1X��dВ��W�-[��M`t��(��7�}VX�27�;ЭQ�.��yM�]*��I%������؎��6n~;}����T!�f讣	В���$%�{B�r�I��븵S������8��y���������gbI$��ʳ��ߵ���"%P=;]17�����~�U��l�����@���&Z�V�XY�W�p�M�~���ٓW�n&B��G��Gp�"v�(��޽�WO
kS4�I�v�!�eR�`'�������*+;���~0L���������(� �e�T9�A$����C0��LZW���\���e8�ۤ�'sF�<�Z��H�O:�������o.��t,�5R���W�����.��0f襺6�@���VnB���KG1F_���h�#k��u�:��Q�n�����.��B���𖂠�2�����H�r�*�����X�����j���-�Z�Tt�e
ߤL�P��&�QD p�����:>�q};��)q`���r��~T����qR��O�`�
����<`������Ɨ��E�]�Uxg��=�ba�����C���<�����x`�isL@���,|�o�V��K�8E6+����%�i�7�����j�y9wt� ��@��L*���!�5�[8#
u:J�-����U\�(����!��}��=����}�������>��,���{��B|~8|8����%�EO�Ys�.�w����"\���wH{W=tA�r`��b�K*ǆ��b{9��	/����L�a��|s�h;���@7�	;6~Æ `~�.7�ӸX-�vBj/�6�� xӟ�$���;w�L�ߙ����Β�3�^��Ym�����j51�Pg�jd���e|$#V%���}�������p�>��/���K�!\	��4E�^�>�m	���jg<e�A=�R���=�Z��9�`(�]�̺	>i���|�i.�J]��g�&k4�~5��i���y��ID��X�9��a�@�x{�h_�c֕[vE�h�<�����DsPF���=�D����ᇗ�Q�G��p� ն����=�����;K9f�8AZ��6v��8 ��:�9�E��$|���_N0:���.ږ�]+Ⳃ9�j9�3Kk}qơ��U)��E/�R�h�/� O����~�����7-<�`�P"g�O\W�غJ�z�6��6;�`��Bg���'��i�-`I4����Ii�B��qS��� )(�M��`HI�O����;��'���S^���(\^��
[���HK�(��h^a��T���Za�t�<��ϓQ�y���JF����$�/�J���ź��N��Х��Z䚝
�����Hỳ]�r�w�Ufk�=?`�7�`^q��ۡ���ID�W�0Qx:��./8��t(K�MT��	7�2W�x5�W�+�[��.�,�Oy+9�a���;���M���F��O��<㈹'Nl�� �բ���o�R����&�4E�@���(ì�F���Y;:\׌0��]��}y.��6�`�h�y�^�EXݎb��.c*S�����:}��N?�4�K0p���L��a1�$#l�����A� &�-�64�{�1.�6Y�Ӑ8(J�H��2<���5O����&%���G�3�E��	�1(�hɦ���C"�oj]�.�M����u�a(Y��5�b��7�2ီJC��t�7jzh�R�x�R�t�Y��r2�\\yd���y/Q<���juAM"a&,^9^�'����g]����3�m���8�V*]�:b%剖	��<�@�7�ɘ����J �%?y/ބ�-�v{�f]���Q��'&�~f��\�T�-X�4�C���A���@�۷y�H�O$�k���Qv���`���(�����Ƙ�@���hzZ�>Z�f�2�aj˕��/¸R���
W!#����#I�5J,
č� ����h��l��w�5�.���6��W�uav�Dp���4��3"@�ݞ��S"�T�ꢥ�ZPY9Sŏy"�$%�E����ǣ.�X^f��y.aYF���B�����9�ǟ�]�ⲏ�P�j���\�hȮ>�ķn��_> A�D%k����Ʃ�1���!����ej����a'rYH��A�/-"k���XA
@�r�q`���sظ��m��������"��L�c��,�T]�m.A ��t{6�`m��{����i6	���a"�)JF�����:dr���s���
��f���O0�R����t>0�As��Ġ���.	>͋X_�fK�0Y�K��v�Q[Oݧ�d~񀎙ǖ;X}���=fs��������ﲴd�㷇�=BqR�@��-7���K�I�.��V|�u<@����iw��iK 6�d���bW�$G6j���q��@�סbY� (�$�4�`�V�i�r��T6�ZF�O�K�I��YU����0�)�O��x�fu��oV�n�P�Ü,�Y�[[l-�����-VH�	rF�v|q	Q�.=���$䅞�I�|����h�������=�gf�����
�	�
���BP�oqVƎ�|���*�$�n�ݯ���.�N!�4�9��G���/�s�YG�?���,J�[��1Ӥ)�Da�W��Y��<7���u� #`y���$�ඳ�"%.�rهړ��|�Z܎�a���چo�7H������~T��ze6 �9<ЧǷz�������������Ӏ��g�¡G�����m�����H�$qY���9=8��E·�]hh`�f��O��KK*UV6����}} �v��
+���ߴ'R�C|36�SlJ�H+;�g(˿�nxDSU���L?�I~����o�x����0��{8�"��(f��'=d�jV���gl��Ѭ���Z�jf�%
��� �,��$�e���R��z�oOP��^������b�<��*�#���­rE�C�}����Q�9V�ԋ"a�᳭QX�$V����&"5�Q��2�De��7E2��&u����2��
��O�~��^CN+bT���K$᜽:b�*�5��������Y�Z�f��Էv(4 ��O����>���Yܠ0�]o@�}����8�s#@�/g٫r&�*ک�/�@Qg�a���%Q��p��=x�y{���}���<V#-x��~�)F��G9��p�����@�sj��AC��(���I[��l0g�(��_�	��-�%�M�����xO]�%㕪�yz~���s�W�
���w����B Y�N���a��,���}|&������^��f�k���	d�����!E�RQ��Q[��ztf�d�m�j-8kc��Љr^���k��]����nwtu}wY�����<5����e��i��%�G���Q�!�֧����`p.��c@?���z��?�_��v��r�r��R���i
ȍ�ͪ�c�n�O1�Ӊ��������Kg��D�!���;pFV�Mw�����_�n�5���fO~�yq<�y� yv��{��V�	�?l��#՗٭���u�����>���-�ܝ�)��V[�J��hb���f-�ٗd�m	P�Pv0)�Q
��������O�v�*�����Ǹ��z��� ��a{F�)�����e�Ĉ׆F~���8!�����y���չɊ6z[�J ��?��Q4��E޽��K�F���xk��Ƽ�?؉x�&S�F@�d7fXo�%��di\g������Gz2չ�͕\+|?��>�F���`�����ΜSYa�s�F�"�2��)���}U0@���6γ5YW���Yv�H���~����S�UT�Xhp��/���tcFh{�H��'f��	������b����|2Ȁ�c�/��D��1�o鴖{x�dp�(X�9��~_f���g�r�#�plER�~Z��#Iq�B,��Z�����t���|뻑�FJ}Щ:4���>��f�~�L�D�5M���ǼiP;�̬�O��,|����v��e�
7�@�*�-�&���?��_�qBv����L��F@�	N�cUfb�d��dK7l�H�P�&C��3���q>c(�`�j��s_�]Q�7�6Wc��M�&[���q>��<"�:���?�n�ʃ��\���氨�v�@q@H�g�{:7�x\v�?���MOq�l�[�y��s"���b�T&�̭�L�w�m0+I��Z��&�_�����Mۙ�kn�ҝ7���A�GX� ��>xqEW�b��I�-J	Z�b@�7��; �܉#��}~%*���BL���-�mB_�L䨛br��6����nZx킃���Gu�(ԧe���-�<�1\n��X��p%G/RMH��9-�08��F�^KC�
-O��؇�q+JW�_�4V�+�"�An婏��{T/��:y�<2<�n@<��#W�g3m���������	�b7|.��C�{� 1��-+n�_�E�Pq��G��)v�D*t�Rt�q:G/��Sf�Q,_����wy7/���C^
8�	tFm��'s-�"�`f�=����z��z@�� �B8$eo�5ŀ�6����K�2l�y��'��� ͿN�(!��@�o�B�z�����W����V��	Ds?�j��ݪ@�4���&�;�0����t�!���d�������ۢ�8�>^x+0�-A�!�b�#r��B��u�c=�!�^:>�HG�4_�2F  ��gGh��g%��XdnL44Y%A�b~��	t���v��C�*�8Y2����dYW���?Q0�nh^����y=��J�o�'��Y�z���c[�O�d!g�#�{������kF �j;��T�MX� {���{���g%����I>Y�up15s�qS�9OY���Ȑ4K�S��T>P��^�;���.]��
�v�Op�^{�>�ՙ{��<�^��z�c�D*Y�攅�D���1�c7�+@��@���cU<1��m��!i�Ako��M�V( �t~����h�!ӛ�d�ף>���m������g߆$�U��ץ�Qǳ�Q���X!S����Z̙K}���{��8�b���G��&ڒ_���R����ϥ�Y4�lR˗0=G��C��p�\LK��X����;N��D���4��9|�|o���'+ԝv�y}���/[� z�n���CΒ�%h�`Kљ�`
Ǆł�^�ߕT�n(�H\Z�&\�cQ�a�e�/�'��|�=�üy�;N!������Bn�h�TJx�ƶN�����U��v�Į�btP�Գ6�U��z�ѐQ����?��*Z�l��n�-`Ip.���y%��\�>J���a ��]�u��:p{� 5a���v\��Z�R�p'�}���|�J�tK��2K�N��a��\�G����;
��/���3Gۧ��"�y�2	�Syxo~��̈́���vi}�8Ĵ���9�ef;���W!*!~l�fI����ӑ�q ?l�ţ{#��$�G�MW� >�_Y�(N_�X�8Hd��$����#a�������rdwn��|�E!� H�������
g|�K�o��,0i.��H�;ɲ_����o�X+ ��0�Ia��vK"�./꯳VJ�
f�=K<]Ǌ�(�(5`]��C\�0�.[��_3��mM'X$�ֈ��VF<��!l;�d���v��R>�g��'O�¾�f�A=�<�٥�M�+\#H��`��3�s��f�SW��ؠwS-pA�-Δ[i�݆�m����^ov�e<��)��l�n�.�Ff�\/�e�����i�6�N6�,QU��ǿ/����c�+nr g�j�q��)YU���x@��f��K�mA+挨*� �����z
�#j6�����DmUD��<fܠ�=5V�YZ�;ҁ2q9U�@]l)���28��6WpZ�H�x��p�_�RN3�GI@k��~�P����L|�5Ê���)dѤ�b�̐�M�,"�Y���mym��#j�[��5טz�6��u̐�0;!�3Je���=n��qD�H����7|��O�MfLO���[fY�Q�no<��b@�dm��O�.&;�o����>�ܤ�E7�ܝ�ݼhn�G�]�P�Srζ1r],��:"<�%�=��B�������5��q��;i�ž�L� F��gG(���8�V:��_�FP�(Z�b�	6����\���N�q�s��"z�T���5��M"\+�%a��B����+�}潍�Cጅy��G��� DO��t?��[�E����2��U��W�z���m�Ȫv{���F<��C��o���Ac��<S�
#J#��3lU@_����De?ɉ3�Z� Yֶ�q,��H��S��;�,7�%㣇��[�2�n�"|����xa�(���B�̂�,q�Q�S��x���c��l`{,x��ć��(u�h��6mpoa��3�7ɲ����m��\c��paC�v���t�@��t18��b��de�0ڞ1xpݼ�a%C6��8�!9J�ky��s��e�8����#Rx����|�|T.�$z�p�h��p!O�t>)���'?VB��y�>��9�{-ձ��������+!qr����鶞���[�+�,zk�+ �9��q���`��cݞ�}9���?�����_-�?t��V
#�Q �՟|S���hdS6��^uo^gr^�oI>tD�����Z'������F.��6
w��b�㌘�X^��I���~h5����^l�I@����(�������?�1�c{�EoN;׷�А��4��i0��=������d�[KL��
&P1����#|��3��SB�t�����餗kL�R�>��` ���1�XfS!�_u�d.Z��/��>��ڄ���8�N?�ʨ-N�z�y�!,^��$V���e�n=叝`��\�XH�#��Ūo�7�E,�V�̴�zoD�:Z��G��{c�MG9���:�L�q��a�l�Y"��e\�k���o�&N�@�i`��Uy莯�R}�i��ԇoT��<y^�a�qkGD�=q�+�����82�J�XO�5ZVq><j���z6	�HQJ�gv�&��ˌ\����#�S2����y��l�:ˠ�W{�t�p �&�R�^Y��k��#߄�e"�W�z {�J*g�">c�q����K���k�F�3͐�M��[>���s���p	�?}F�N�'�P5��D�:�TQ���ڋ��.�4)�&%xn]F����ч3��
Cy���5�@ؕeBX�I���ʻm�9%���h�:K(r�G�I���.ܲ)�Գ���v��ñh+��UD�_V'��7Q �\���)��?1eS٦���ZA�:�X��g��0�sE�tn���2)Z\(D���j��H۰��?v�I���0rY��F�u+�-s��ڸC��T�`�,�Sx�l�����̼s��^��z�O����� r�qC�FY"h�5�/�L�PWfO �/Y��o>2��
*�hFv�[��5(�S��+0-#��{P��Wr�OAX���A�.�[O�2�W舜�l�fZ�bڢ�`���Je���l�	YVD�x��)�nf�L�F�Ё*�ol�X_4�zRw��N��)ĥ$���g����⹻ ��#��~H1D,�M�1ő�A��<#��uc�7�y=u�A/Mt`���M�?Q����J��t]�|g��!�Kc�:�.�T ���2`�-j8�b#�q�������
�0u&��cV[�{����R"�w����5���T��������T�� �[�2�y�ԧn���'O��DX� _d�mcw�~����ݿ�1��v���h�
��2�b�C����09ˋ6i�h+_IЃ�|�s�${�vN0�>�0T�&��gFb�U5@�)|"w��S���Sc�Ť���i��R��a������{7	��>���z@1�S}�����V91!~������q6�E���6�2������Z�d=̀�Pą����e~��<�i��9�.e�+�6���KE4����<E�4�c�F�e*g*�zϝ_6��6��£�_�jE{��6+�P�X����"���7��&�l�ό)JtF��<H��C���}0��e��&�������N�˛F20��l�U��߉{��]�W�J�B��]���\--�~8�t�������L�	��T��vș	k;,�����z��L�l4�V�.�8h ΥA.O,��̧lN�Y(��^�H����W��DC(T��97��=��f�:��kU�UL�Ru_H�����ُ�cu��_�r3M^�uJ��v��!�	�I��ѩi;0Ax�=W�[��h�`�s�S�Ѷe?�p�Rv}%L���J A��=@��+��z����$��!�lV�Y���℠{�|2�W���Xng�k<)|U�SZ��꘬�J������q8�` f�σv���š��4�j'�*,�,�ʧ�ݙg�Ag���UHn�j⟭�t�꼂�!�+�ꐔK�j���3nq�I��V!Av�"aj�&D`˩o&�	�e�y2��OP�9��Ezr����i�[m�s[N�焮oF�j*p@/ �e�0�ky�gD8��8�Kj-�ɬ��U�~�j/	w_�VWb����\;�e�<�%����׹/����1��Ls3��a�'�yE��1&=[ڦ(�����fd(��+տ]�k:�	�ї0f�1���篬a����,9���*�(�z�-%��0bp���זu6%xd4$�V��"��PB_�ܳ����N�,\'d�	��vkX˻�0('�;��=��y�k^������T�V���C�Y90�f�qn�V�2�5T�b�lgt�ϒD���c���t"�����X�-Gst�b�:L�VH�ib9��ցnvŕ#&q�mim���
��b�� ���E�p�깢D��"���w�1i�U!��/ks]�?kє��_�-n��?�����sJUN��,���B�����u+��D�'s4ՙ�WQa�h>����ۅY�n��=�7�)-�@n�<�l�ts@dV����݅�����g�X�h�#ax���6���}�B�Ba.�}1ԬH�vi�S�@�B�S際ᆵ5�6��kრH��&�:�b�MfUTh�zAHF�s�Q�Al�t���&a"+zh��,�Q�:P��^�3�7e�\�E	)�f�I����ȯR(�@��`��.gT�Fb_j��).��GZ��X�
�t���? �����e;bq�����\����F�Z��/OH���o6V܍�Ժ$�ߐ��
C1c/�S:�a��C��lE�c��������rF�,�]b��4>$/I�����d��ғ�q�)�B����\H�$W�Y��nQŻ��ʥ�ʭǸ���h��p��l ��r�
{ 5��b5�E����M�|�Y#YZ����%|�7v��(ҀW��I��}�2�#$��]�b7�&�Gm���;=!B������+f[Cmh��
J�Pwu�V�cX��ξ�+3"?�,X��s)�-�c*����@�cst��_xH-~�<�l>�D2\�����io���5F�V+�mT�k��b��e�����	�Ȗ���S|��>O��������ۀ}v(�5����Kh�D�i���Sr>Ѓ Z�6[}S����++��Q�ڲ�Nܲ���&�7�W/7�����/4f�fZ)M��^�Ɛh���V�ڠ����V�h�M�ӎ4��ך�MaR"�P��$���3vj�=Ay��ʝ ���U�8��{FG���U�l���I'v&�`�eO�\�e��z�,}�[�j��>�k���0���/����	@�avO�����7ӗ�rټ�1����$��8�?����e�����GN��XN|�
�f �A~ �զG^���k?a�ȎJ�C����|s�y�����������;s`�H��3��g�jA�����܆۳@T77�Fw!,���㒀"\���&�:�Cߨi�g(��HZ�(?O�-�M�ú��kp<��q���˖�Y�*�͆0�>��qϼ�8��t05Y�I�����3����"8�]K�]롗�8�DJ�u�>q��V��9�&�i	��·�Te���P�ˇ+��Q�{?�h�[yY���逗�h�qg���z�fjE��fД�Y~�|/�{)w�mVĳ���9�Zu+�R�о�t�Zyϩ)��E�L�J�ު%ԣ�Ւ\�?�zg���@�m|��C�=����y:XV_R���]ҿ�.#w��|��A/�%a���D2P5	�soږf'�v"Tz���b�i�qT�"<AI{"SṇEV?+��x.����)f*���qr��f�'��'�}� ��	��.���l�O��m�d�MR��
¦��}[_��u��>jR�
Cem�:��ש?�mOVԻQ��rl�C� _��K��Ļ	<���U~�	���_ػ%��u�A
ǁĄ�E��4��3��������x/��t�q�������N���j/��f����ֆ��5KJ+M�_��w O��[�R��P����L�;���ȍNr8�*��}ċ��Xܝ$�U�>aB�\���֑��S�����$iY!�h��2>��&Q���c�S�)6S�@רl�"Q��8����1�<�1��k��yt�SO�n�{'��BVe�{?��d�R�A"E"�Ӥ�[��x�ݝ�G2^]λ܆3�H����
&���B�&��c8���~��c�-|D�݅�ĸP^�b/ݬ��쬋��o|�_�E��i����{ �빂#S�mX9kJU=w��_��v��C�6K�]��@�=R�æ�������׍1F�H��D�A�8f
O[�G�'���I�!өqݛ�U�l�u�E��,8��2��s���{邹��U��23-
�,[ĵ	vf�i�"\��W-L]�	�i��ʃZ*[��������&{
��ʭ�W�%�~.�X��Wu |dĄF�Q�D�J#V#��5���k �q4���:�y�w�Z����l�+���갭D|A&7�xg����Qh�����&3=�`�x*�B����#��74�������3�0r��M�15�������F�������*Z�ǁ�HM���u��TMj�>P�1G-���]�� �������O��������  �ǌ|~�����@e�yN������6�����,<w1&�<h���N�aat�K���8�ҒF2�>R���&��Z�нh�$c���Hs�Ђ�\BH�)��|�W�4%���?���ca�$�H>�A�
�,(���mh���V��<�x.��'�����*��z	���kt��n_����S6 ��$m���Ew��[H��=?��'�mj_J���)��;�c"�Zim�B��%����D�J�����j�$7z��H�r�S1g�[�ȡ�^Fl|�>/Tik�Nt�r��#I��UVG��o9��%�T��Z Z)H4W����cA��Rl)pha�Y�Q��IL�'; y��'����$gt�
�0p)�_�^��X�}f��U�˺���gɌd�P���=˾�4�K�E(.�z4-f��Ѵ['�o���y	M)��8�Վ�ęV;�O*�m�~y�zSၦ)�����k�>�W��}��{�MTo�^���u|��^�,�)0#�r���=2�c��w���;QP4��g43mc��-����#>6Ҿ�x���P�8�Z'�[��
�!��A8�9���<wV�"h����i��W��E����M߲k��8I#�n`���iV}��� ��0'S{�R2o��,f/0�>��c�NC�x���S�I�:��W�� ���G�/��U�����$��,Y/?�]�Y�rL���OMO�������WԎ��E��������5����`Ē�LC.-Ć貧�p�P-�}ҩ�]�)���w����]�0!B�:m���B�A[�k[$)�=���p]�a}�h��{�8�,^ո*��R��3ɶ�z�ǿ=�Q�t�}�ʛX�3�������6��s%�������?��br�~M���ǡ�|2�m�!Ϡ)`f�I�8뜚%&��V7)[�����p5&zy��@28��.� ��X���$iGY�mb��.���̾�PQ�5�|�ͱ|p�iO-�}�[]-*�^�%�%�p�R�4�	��.�6DU7ꀘD��
�@I�j����5� c0Ɩ�������"� �B�a�ɧ'#�f�)��(�o-��4��dW&)���v̫|b�:��q�jX.�����Nߖ~) ��)����O�TL"�1�V}D:�AMпZ��D�W�ϞU1&	��0�R��``K)`{�Jڦ+352��q�µ��	�E�x���u��O��3�Թ�I�,�b��F1c_c�c�RhZrf5fU��!s:kJ�7�0ɯ+NWGG�Q�DM��e�lCX/�m�=�?C�I�V۩��u� �� -�4������ݽ޲?h��աL�!�o���$]Y:�Y���7��7f�KZW�}?���n�TT'���Iՠ����Wã��#RO/�K��T:+y�Q1�5VkЗ��2���ἃ�N#���� r"ҁ�8}�FmL����`�Gdu�U���ZIl�N��+2
. (U���2���ǆ�r-���v�[n�p�$W+w��b�wy�W�[�.�j���hv2��[ː�ܼa���o�Kk�DTv���P�7B��QO�ں6�{�̸�lU��e�����ⱶ�s�5��<.��13��(�26X���9ӳ�|�VD�]������]���������'�ȼ��4�ބ�	*�lQf���c�ˈ���~��Ϳ1g�������J(oVk/lt��í!6�l�gg�����=�C��d�k���>SDN��s�RY����P㏑?�0t����n��+)!;�T�x��	6�������%��f���|rG�Ƙ[����� ki��zF�����t��O+dD�[���\WM��O�8����I�����-���8e����(�B��O�5��гu�ռ;҉��D���x��\��k�Q�J:�V]g���6�IA�d��o	��-wn���M�F���N6^��_B��&�gN��oBx%���ԍ~�1����%���w�?�.�BG�(Z!�YsV�����,u�H�.���]��2�N7� <�X�Tx��E�v��'\|C�ǈ!��G�c{O��,~�+lpDT�6#1��"�(o��z��>��!ls�)	�Tz1՝2y��0��M�O%5(��pL�� 봋r��W�����lBve;-|"�]�狅��/����3;^�Yó�\ْ�ٮ��a����|A.���	��[O���x��1f G3T�O�E*�鋊@g�]��ǐ�{a�3,1_ �lL�͋�UO��C�uiH��-ƓXtz�â+[	�A�=�<���'��I��j��0�u �}<%]j�9_�8��~���Ba�5������^�b^�Y�3I7�����B4��v�HʘT�gSM^Z��*c�3�er^8 s��)�
<cm��o�jE���`�&��@��.5/����>�5�qbj���:�8`��-�V	��_̼�������k�kw ���sG����7��-�	��{�N�%W�tH�CE�4��e��Qv�(biji#�8n.�T(�)��h��t�3�}�]���(u�����Ԧw�|7FG??Fꈹ��2.�z��F��ij'Sf�%��">���i)Vך�eע�B�7`	ƪ'#�_��%��O}r����ǟ����{��̺�L-Ф��{e�4�Q�\T�AA��Ru`m�}k^kPI�n�&�v�䨞u��g�/��Z\\a�y�L�$�j,���RN�2��0��&�G�G��E�c#q�7�g����N-YUI]?�]�r>~QS��仧�]C�2ɥ���s�ˬ�K<��(��[@�n.��f�LM(��j���7��������Z�[��|�q0	S���X(#>P��'�L���O�G��w_z��+5�����5J��gGP��x�4a��!�U��`�Ի%+��*qQ�,Q�=�}�q�S�\.�iT\$��	S����O�J��<�,Ǫ���	����O�@������[h#K܏c�j�9��a	w/,\`��?n�
|t�c^|��?0lK4���|C1['�'�5v_��w���Ha��HyB�*D5�BD�-n�M	�(Ȍ! ��
�qޅ�-�V�ȕ$շ������߿�گmI����Rl����k������o'dHm;N��zĶ��A�-��H��^e$�F$Z�ª	y�P���xy��M�:6;�9wo]���D��WO|�S��7�J��L�hU`����=S�?�(9+-���ݯ���!d��{n�;S�-{�!"&���=?��嵡��4���L-(�G��5���]/p�7=��G/3�S�o�t�q�7�������c����9��c|�Kp���&`ɒ�^29n*'�n�c,���%�$?�!c�c4�/*fr��\�Gxǖ�*��q^3wb�uݹ����7�@	;�F�vE@�[�o�,����J�8������f�i{n3�OI|�w$sC��I	q��wS�PXi0-S՛�d���B�����]�'%��9����ss�Һ�w9����\$�7�a����_K8��jM��Fg�_'�h�:�H��U�#�z!H��1���Jdd�B/��L�����~��DtfsF�DL���4����r/]:CS�[��N>�C���¹�w��p�8�%�ӷ~2�KcK�_?}>Dl3;c�w�~荢\��ɕ�Q$w	 ��~H�MO�e�ɯ_
� 
������R�h���ozB����XB�ʟѮR�����$|"�o%�q�9��;*����hv:�S$������H�qO([[`em+J���^������-\�I��J6���R,8]��qN��L4����m�X��bץ��B�j��=�P�f|ꦎ�)L�nk��	��p"��x�:ч2��
�F�_����m�(��u�m�N W�_��O=����A�{<�a	���m !��Ν���p�	��g�n�g�s8��Ð�J	X�=F#P:1U�,ݭ��Ď�b^�[ѸՎV�AS��Ծ��֟������W;������ݘ(���oEz6�;��&C���Y�y:��sNM��1<� ӓ{�y��������P>��D=�\H@s��~��q_���eZ]}�_���-3�һ���s�vɮ�eH� ʏ�a�H��؁J��g�#�eW"r��N��4��g=���v���}mn�b�]�g���X׬���Lrj�Avp��c�o�tFR5.q�N'1�s˧�T��#��unBU�|j�d%�:0=��/�~�OF���b�P�C���<��� -:9�Py|�L<���1�AB|�����t��c2��M6Vx�c��<|R�tU���;n#����q�Oib������}��-4�:��k;��u�"��-��&B���x́���9�Rݚ0���~���	���A��v>/T�&݈�@��Z���N4%��X� � |�)"
Ek�6dz}R��_�{�����W�Q�PrC�^��6#��R��e���縫�� bq��-v���i�X��#�����4�)e��REu��zF&>[�A��Ji�=˷����`�,�Q���}���f|���G��)Xȧe�i�v�Z����am��=WΥ�����b`_fU��WOD�"(~D5M��g1�{"ȉ�F���fxNF�Q���&�}hہ��Aq`�
����	L�	�>��x�6F#�$Hq6La�a�R	�&-G&ǊoYݺ��n^����gA��c~���H�B���h*'�Ԅ�p��1�fJj\�"h��Y �=��	Sl4�e�E��.��X �o�;#�c�@����Yߎ2�/��[�fTk��ԩ"=��/IruEotV`F|#	MȾ��j3C �͌��W��__�u�Z~����G���iF��WD,��Cº\Z�9=j]��m��ݧ�&^��A�/�#	��q�_k�MB��S�u/o<Ӛ�}T�Y�_ ׌�f�8m�d��(��y�~��:܋�e�4]�{�Z;�n���Z|��0].�}j]w���QW�Y��F5H���4|\8��r��0h-q@� ��`\8ars��/�q�իF#��U㔘d���k��	���iX��?�!���λ��[jh7�-�tO����n��������qY�����wS�zE/TŻF�A5��vz���}V�C�c'�*�*aQ~]��W���{$����ڣ�H�|��{J�y/L<��y{�Н��ۦ�|"dAy��uƮ������1�00����7*��ۚ�ּ䟟~֟��bi�6�#׺�
�S��h�^��ګ�gT����W�.��t�bY�E�[�Ѭ8������t�H`������:F�m�.%������֜l4����n-F7���� ��g�Se��4�܄����SI�#.��kP�\LIp�g=��k.4,�,���Ot���������v��{�f�jc6����v����M�6ޏlIy:�>��e�P��ai���z$��p�@rQ9�a�-�6��PƓ�z�mDn�E�vɄ�v��@Tqe�~�cQ�������,�L^J����S���� �{�'�ޖ�W?���v���	B�vΏd���9/�덬�����@t��%��\�Q� i��b����D��b���X��X���Q�@����)���0(���ս��Ø4��4^��O�lT�G��iގb�5�o�������xJC�goa�(4����X�M�]�u�0*�O#�)�;��B�ٱj��{�PLǀ_�Le;����/'~�@��Ԭ`�o�`&��=��Lک/<�bfحm�ؠ0��O�:RM��&rQ19���SU��LnWX�:��3��h.���u" ��I��:�}����ѷrf����1A��ATJ�b�1hz��GK�~�1��V��!R�ĈX^��h+��	�#_$��`+��Y��b9#�b�`�6�����£L��k��s��}M�{��H�W�ͺS8�:nX�������������X�}>��k[�w�Y]�֌p�p�Jgp�vY�E��f��
�g[�E�������j��/A��#B9_.b��.��H@kZ�������LTD���z���n�,	QveV-��6������_h�E�=E؇ h��)Q%aX��L*��/o��,��۠lk
�	QW���%�+ڻR@@�+B/~�WѠ��g��5E��:Wp�����Xk�8u�a�&k6��O�16�{0X�Aۦ�d3��V#�s�@�EY��9O��\q�S�p��d�k��=[���U?sQ�lb�'����ERJg����Ic�@S���o������E����s��n_���yl��+^��5O�NZ}6�_��5_Cle�!mH���Z픉rd� p~
��=�l���rEs##mz��1θH��l�	C�VD6w~g��b�aa�LGk�u#�g�ß�����+�..2O��JUH�{�w���XD[�s0j�1P��e�(?�i�Nʓ�%8��������VjdA���C�^����#a�̷�)�L����u��bEg-����������w{�Q�a���Av�ܴmR�	Rb+T��JdukT@x*'��Uip8�SʱZ��2�̣D�R� ԰u��C@�m�cK=��fi��ID2bې��;�l�����G�Qnp���𼉞�x�E��?��>Y�Hf��7)_������0ʳϴ���"}[�����GNx���0vAaR
��6
��u5	$70�D��b�h�a��'(I
5�FmD���
P����P��d_^�K�	"e���F�H�u#.}�e���
�*H���hU@�������^&����ȀBε�%ȅ�`1OxAQqP��������7LT������#�1U��GM��U~O�[fpe;7w278�N�,��j�͒�{�NPab�X�oԌ-���#����gs���J��CQ�y/.M���k*�Dˬ�%��l��6{ً(���<��x��po��*�1�.)$L�Y	TM���Bq,���Mh�D���R����M���?DI<
MY�
/��у�Mx��]s���|��Q��<��N�M�Y�o�wa��!�
�f̟+>�@'<�F�<g�L��2�ݱ�,M����23Q#d���3{����8%�U���d��m����+�c�~b{���C��XԜ&��EVo�H�Q:��QG�P�R>|>���o�0X^����U��Q3��Y'\�&kj�t��=&����f��QT{��8I�se�w	j2�n�7eN�6چ������-Hk��s��H�j�J������ǜ��o��ár�����d�4�a�ACLr�b(�k�70�S��Oݴ3��H^
�x��G4`Jg��*\ܽA������N�&�=�}K���
d`ֺ/SE���B9#��E��?������M����\�3��z�����l�1����cK)1��^�C81榨�`��xmo��D�U�Z�ї�T4��Q:�RОs ���ms�.�V2�������1�w^���p�\�%g{`�w�1�q�� f����G��9�r׽8`0&�L�G�$�mBz���o��Q �B��Ȯ�J�Vp������(,�
_je�:j�vZ�L�`CG�P쿐�	M!�3�`�wѷ�����7��_�M�%�l��I@9�s��΀�AɗY��|��Ş����@�`�r.oW8]�g��w�ބ����wM�	u���W��տB���S��B	h�?T�^� �(���ҏy�?4\&A�i��|�H��4~V`�� ��f���JmqR#���ʼ=Z��2X�1l6��ƿ7��O�Ӂ��%�Y�{�̜l��ny"[x4f���0����n|�	�4BB6��KUo�P�V���Х�4.5�ӳ�(�C.� ƛid�5e����V��W��;�`�'�&��Zo�B��W��đr�u�j� �]jǛ��E���Q_�UsCʖ}y�����yD80�V�%�>��ip
�U='��O����]��V���Cr�1���H֎��Ei��g�w��W�	�د4�?V�Êg�wTP����������Rנ��i�U��z�f,�<s\�:��d{4��_P�N��Jv�6Xg��e���PRz-A�=�ʢd]⣠����E�r�,�ͳDP��bXtf6N�aT@�5T�Ao8!��6m���jqA���3�W�]
���f����i����u�h1ş��I2Q]���K�8�����L��V�p���鄁��b�)2m��c։q���o��Gk�zǇO�Q7�ל�r��*T,�p� �>��q@����Sq
����2���7�o��}�Y/O'2�Xj�����Dj�D�K(��ZC�q\�|�
�=�4�7�V*�T��g�k͏t,�H���KQ���	���yD4PD���9LC���,tD�ǩ��]An�$tr�-�H�UB�h�;0\N���/3�b֢[>Cw�E�w���xR$��0�8,~�t�Z�0ͺ�,���]W�S'�x�ßnP�Y�is��Y�����Z����Jx�}#p��Z�S��{;�-UG|���ө���)'���������B=���y�=���v'�V���o�L�zR�Ղ�J�h�/��Q�3.]�
���O���(��
�|�/��!���4*ث���2j���S5��m��` �f"��;��\й&��vl�S5P'�Ad�̎���i��W3OE������R�Ĩ.�W���G���"�1!6�q����*�hr�L��U�;�8GI!l��o<�8��
�����UC�l���r�M�Q��͒f^3��R��͔��b$���q3%�+��Y���e�_4�<0���Bo��_N�!��za��<��_6��8q�³%���} �t+��̍��Ek�"�ִ]�(�;�;�d�f�ޜ7��Rz��]���8%0lb&6�|ƫ���[G{VV�h��Ný�ב(�o���zǳU�)��X��!���������9��������+G��)M��$��q�U��KK�z���8���F�TXJ8��K����YWW�3O��9bj	���mh����Z��xs{��{�i)�����}�f �(H��͞&�b�{����s5n�4�9�)>2/��@�U��w��b U>�|h�?�@�������HZ�[k@�V>��/C�Ȃs�m����hm���⟔O�=l�g��T��GL1�`���]D��;�o�E�ao_�� �xPK�U�����b�ō�<^a�����̗? �_T�=_��#-|�/*��"�Zv9��5�eK(Z��*>DL���Kk��Gz2e�s��9ua��~|��շ��Tl�Ɵ��N�;��=[8����. ��a����l%.�^����U�d:�eߤ�*���#��J��Ɯ̜bb����5R�h���]���j𗬕m�Oρ[�hWr,򹘦K!nĳ��t�*��p�X�E`Pg������^�DM�
\*�ȑ�ǉ$٢#"b��|��M&�v�?��WYj�~��� �q�9b��#��?��S�L#���s
�-O���%z5�k΂r�I�d��P]6�в3
��,�=���Q/�C�}�:R����ׇ��cZ�.8��M������+7ܒ��te6=Η�QS�f�0�zd[\ݷ��S��j$M�.��I�!a[��j��8�"��\�+�PP������mu���acn��Zv#"W�@;{�������^��e��cUT��5,��y1�m�(O�q�bvw)�ѿ{�W//�9-T��#�D+q���a{Z�5�C>��}١�۱�"�WrGkz���{Ev��p�k������7}x�\�x
�i��V*4a�%�:�rr����&�]������(�j�өՠY�#C+ӽ�Ů-��2F=��~�Aٲ�P����ڇ̵� ����beMa���w�1��|�1^�N�޺�7�N��y���/�7H���߀5ޱ�D8���bGt'�a0�@K���w>ZyJ�2��]�7|��Q4�1	U��1qL7Ӝzټ�>u��+�۬}ͱ�,��$$r�~����n���c������R��������9�Aw�WNF\ߨ��	æ�}��>����=�^�D�ԒlY�R�&V�?�+#�r%��4�A�5���x@?�������	�f[�K���m�5ܭ1��3pG���n�(�%7���`��iqt����,ج�^�K��8�`�u��̀���0=B�3:b*�ib%�~i쨰�0�tc�?7v]�W�wD^T�wT3o�Vz��$�	�l�m��x=H��c�]K4�<�|�
���{7��/p�-6��)f-[R�w�O;�y@�m��q���N #Ӗ��̸������_�����]Y ;
�3����1H�!���`�광��%��LD�ZӒN�Ay4�Mk�b;��Z�&I���!��i���T�<�A��JoH��î��~����G�{t��9xD�X�Ͻ1쫨q@g	���7�8�%F��nv
J�XB-" x�S�%�������a�fn�X�$���J��G���[��
����	>�h4`\x���v��@q]~:2��E&v�٠0�F/d�mא�̌�����B��U�1�C��by�Y��,���Ĩ��㕒q*�Ė4�J�z�,�u�`���Ģ����5��E�� �U�'���J��7#r�#����W�ߦ���fK��sF	U&?�_�u8g)�C��h8�X�E|�>!�$-�	�m#��
/����'ڮ��Ł�|�q'���[�������X���T��������w�M��%�k87t���S�jI���*�	��Oo;�Z�v<�	��og1=��-����7�$���⧫%���~�H��.����h�-��c����&MG5v?���s���C�$R�A~~=�K����BK�����*���������`eWo��hD�z���V��e������� d�m1����\�7a w��cK؟��_'@����^MKc�
-7�Wy8�(�F�e��Z !����)�4g�B�������[�{ֱ�/�8b��׭����yj�97��*��qA(B?&��!��[J�ڄ������ӮALKC`	���W��--a��oh}���A�Q�n6�Z߶�� !�X�2+���W�r� *���w��.I�i!&Ğ"V��(f��U�-�1�	�"AK4䊀�JB}.[V`MgJ��JqsE�%��B��J6���|Ǜ>�|�Qoh_�xʱ���tZ����G�=�AK+Ԝ.��b�������)g�Q��j2�y2�hS�&@K�C�a�s�]f�#��k�	���a�������Z����ewm�9���^M��1`I�������<���m��"ϰ�g�|Ҁx��+j��Bhᖋ�RG�Z�$S3@F|����텇���%N����o�m���*���sH����	_'�w)Z�ݯ��0���z��a�+OE�����]w�B�f�9����?�}c-�Yј�)�:ks8����y��nJYᾖ�`cɇ�ܸ�l�Xl��т�［�Z�h%�Es9(H����%��Y,�g��7��:��t�nT��^{S��a'Ы`@z�uʻ�����5$1בL��.��5ӯ��l�d�K��碚�)w9O�58�2�/���\m���ifM���PQ�!�혓�	(Ql��|�e��1  TI�ݱ`W�L����� g^�d�h1��L9͘7�-X]�i1p�lQ]U�Տo����~�C1&�E�GvDy���g;	b*�9ܒNOP!���&V��u��yxFV���AJ�;�DM�m��K�k���	q�e��	˳��F�4��4T����VӀ�T-۷��e���J�����Ks$<��=�p�Y7��w���t��M�w�ވ3_0H��)`�B�K��
Ew� �b$4Gܿ1@�a|l���̪S�R�>�gs�&���<����0��B$IP��&&OJ�e_�Q>A'��ޟW��=��*T�b�7EzYE�o��ea�)I|�I��Z�0@�G�/��ш�G�R+��gCnS�KJg�.��7~�:'S�N�V��kv��F����%����8
m$�Y3R�@SW�檇 5��:��q�3F��㺱�t5ҦB��k��g������E��z><#HT�Wn531_��P1>���tD�[�V���w�{�A�t�r�KJ�$w�(Ci��;Ӣ�p9��!M5F��u8̳d����7�~f/K����!!a�o@�p �}���]��dz����U�lB����nc� l��e��%OǍ��C1��,1&��3����4�^��SZ��{��U:�<��Jv��J��O&AH�����N%��<Q�H��{�F��AWO�a��fW�/F��^����<��q��Kΰ��7��g�V���<.f�it�nQ�c��,����xR���S�P���-Y�G[d���CNC�'@�ѭ��w""�Z�{,���l ��L�C�� '#�ۯ�5�ݓ:@��L�S��.b66=���(��/0=���d��j�W!�G^���f�\�R
xh�n E�qn�g�rI�,�PC��)%���Z�>�D@로���Gx�첗�_���	��_�꺄(H��N�|���+��4B���5
�7AMc[g���3Sb����_?�:�'����k���_)�j�B����>ٺG���_�,&�E��T�6y6#k��3�y�hN� �׉����fn�� �S�+��v0aL��x�S�yY��Ƈ65��}+9�Y�ʹJ��t�X�e���v�'*�,��c�צ�e.�xd"�w%mo0Ө$�4����Ϛ�%�=*�k��0�#�a]��B��=��<�~�$��IW���B!��H��>_#���EBg�ӏL^��"�J�w�Ţ�c�<�v�f"u��ɬ�6��{��k*�� T��J2$�{��N��Ɇs��@��=�3>.�APBč�ږx���g�l��	����8�`L����G-!��� �獞B���6�j�,SL�F@��c�RT�.�5�W4���R����R���N�9�ʥ�qU�ﳐ8V����w�����h+�h�m��;��\!{�2J4����牶�MT�����s:�,MZ�~��S�Sd��5��p�(�c��,��&�d�p���]	~o�2e���E�[�$\=t>u�z�66*��nw�f�~�\3��WPRز	:���_b�L����vh���><�XBEr��1��|-�ґ�>�n6��w	Y�ljE�n��N�HNH�L������B�RC�Rz��d`���.#���i,D�w��0JVsUn�j�إR���y%6��d��qɸ�ߊ���,�b�c���&2VC�W��3[5�Z�����Տ��*L��4qJ�-�zC � 3"��f+��@a��#6�S7L��S�i�"K�T�:=�w������>�J�a�R��!BX-.c�,{�N��;q��(����Km����������w.!���Nj�E%��MIR�Vn��y�z !E�q���E��;��8�mG�С��>�߆� ��82@�:wE���mns����}kFp�G钶B���6�P��s�M2�[c י9�H��f�:I[HVUZ��{#g�$��+���yV�������+�v�8nU�R� �{F͞ ��8�Kr���d󐔖_����&É��вR�֓��`u�`X^q�ӂ��}w�O�Ԉ��;��+o�E�ێ^��K��n�+�*�¢j��-�6�pig]�T;�J�"���	�%y`�Tm#�
I�Q�i� ƚE�% �M�aV��l޸��=�.3oʀnuM7\�Dm�&�E�m��L�ՉT���b}F0�|��!�F�0�r�*��?>�%J��5{-/J-�l0�R��Q��o9��!��Zf�V���YM�\	j���]��h"mwи�B���}���G��t00ˎ/�Ƣs[L��e��"��ͼq�h�.�������%Q��f#W�ꯧ���)�!�h�i��힖��U������7�/��ek|%E�I�H�?�0; ��U4��,͌�uD��N��"r'�t÷��T��h�03�[/uE�
��jv���?����SB�{�x+ܿ��u�t��%���]���1��x�'�__�z��_A�[m<��ƽ�]���*�����O	F`�(	�|^��q�l�����	�lL]��̞��{����~��C�̟��XA�C����L.eљ�g��)��;�C"1�H��M��pϮJMe��k����+'����Jk����}��kL�Y�2iϵ�1?�,
o�o�7�F׃xso��xp��7*>��*ӣE!�Q.̼R&���G[W����`C޾ַM���줾ݥ?�v�4�mw;ڢ���h�Cu�^t���4A7g��wk�q(�l�ȉ����K��(����"���P�@�n�%�K�cRHȵ_��<��b��Ͷ��H9!g8�� �TK-
$�L��>[w�l�̒�?��B:����x�W�)s�����W�V6��&q���P4�?�����Y'���s�����r��܉J�`�itE��y�rۂ�#h��>�A�P�w���ƑI��E�[�#��4g$�es����ca��(a�,D��|fQB�h�r�,=P
ɩ�P7�6��@(��_r�������6�	��b�;S��������ۢ"�{����f��-N��1��U��-<`Tv&�g� � �u:k1�����/�����&�g�9ڧJ#r3�P��@G�E��T�Xu\@��4���Gz���l
�T��FkS���.?��h��G#jM�U�`�{S�L�A�(4e�i��X0u���o��
Cƶ5�����Ф�5z��hp����|{)�DR�ER�TfJ2]��Y�
~m�I�@P�M���}�d�GaJ:�,��M��5��/p0���<�ϴk�o*��\��ӣ��UWlQu�>���b�X���$*�v+T�6��Ť��C';)mTq�4
ɭf��WEy���] �/I�z�<fi� ���F���{SUф��h��	[U[OeƄJc���&X��+g�pI���S*Ylk����u�ZxiF%��9�i�no�5Yq�~���=@h���D�� 2�������f�F��h�������#f�x����85�ޖ^g~r �)�u(K���Q�{[�c�X��!q��H$K��f�qƓ.�5a�8[��.�u(�6^=(�����*@����9�f������OFx�`����`2�k�RB�W�EX���_k���O,��C:4'��gtIۻ���~kcf�霛<+�W��H>I�"?Jf��D�7J�`0�����7+�'��ZB`�����5���5�P��PՊ�I& �tG/�f�ʆ���Q�J��U�����'z�s�}.��3���R�詶g����yj���n?��������g*�<�����.��Eaę���as���Ȗ%�L7��v�J0o��}�Y��ɲ���_���ų�.YC��,�f�d �c>UQm���r�Y_~B^�߱�Z�%L��댁J��͊�\�����;�h�!��_���N	���Q�بm/�[7��?���G_f�s�S�Q>>.��a�d� u�.��8<�Zu>���8�Ӓv��.��VL����V�� �}��v�4?�7�m���/� ����>�Zտ� ^��Z_�>�fe�how�ِy��+��2��BxX�ּinO��o�fv�=dw�q���i�@�Sa<y�y�݅bcֵ�`��K��%�z����K��TG^w�Q�6�}g��tV��R���լ��9�S^�������#�ј�Ў�Hk��nı�^2m�%rP;��	C�����f�?��z��aK~X� G��?�ߏY�V&I �6M뫃Ñ� �rSt��Hb�H{�J�7wXD!��>kBW�+������h��|�(eQ�=N����r�݊�S�[D�=�v��L�3�d�2�����'w�I$��";��P�+WV� ����0����@�+���pc~/��?����Y�q���G�te6�uE�Nor���stlg�D�N ��§�$-����`<&����`x��1�3�g��ہ��z!