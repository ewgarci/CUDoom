// memory256_16_0.v

// Generated using ACDS version 12.1 177 at 2013.04.26.00:10:27

`timescale 1 ps / 1 ps
module memory256_16_0 (
		input  wire         clk,        //          clock.clk
		input  wire         reset_n,    //          reset.reset_n
		input  wire         read,       // avalon_slave_0.read
		input  wire         write,      //               .write
		input  wire         chipselect, //               .chipselect
		input  wire [4:0]   address,    //               .address
		output wire [15:0]  readdata,   //               .readdata
		input  wire [15:0]  writedata,  //               .writedata
		input  wire [9:0]   rdaddress,  //    conduit_end.export
		output wire [255:0] q           //  conduit_end_1.export
	);

	memory256_16 memory256_16_0_inst (
		.clk        (clk),        //          clock.clk
		.reset_n    (reset_n),    //          reset.reset_n
		.read       (read),       // avalon_slave_0.read
		.write      (write),      //               .write
		.chipselect (chipselect), //               .chipselect
		.address    (address),    //               .address
		.readdata   (readdata),   //               .readdata
		.writedata  (writedata),  //               .writedata
		.rdaddress  (rdaddress),  //    conduit_end.export
		.q          (q)           //  conduit_end_1.export
	);

endmodule
