library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity texture_rom is
port(
	clk : in std_logic;
	addr : in unsigned (13 downto 0);
	data : out unsigned (7 downto 0)
);
end texture_rom;


architecture rtl of texture_rom is

type rom_type is array(0 to 16383) of unsigned(7 downto 0);
constant ROM: rom_type := (

--Red Brick texture MSB = 00

x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
x"49",x"c0",x"a0",x"a0",x"a0",x"c0",x"80",x"a0",x"c0",x"80",x"a0",x"a0",x"60",x"25",x"49",x"49",x"c0",x"a0",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"25",
x"49",x"c0",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"80",x"60",x"60",x"25",x"49",x"49",x"c0",x"a0",x"80",x"80",x"a0",x"80",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"a0",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"60",x"60",x"25",
x"49",x"c0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"25",
x"49",x"a0",x"a0",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"80",x"a0",x"80",x"80",x"80",x"a0",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"60",x"80",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"a0",x"80",x"40",x"25",
x"49",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"80",x"60",x"40",x"40",x"25",x"49",x"49",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"80",x"60",x"60",x"a0",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"25",
x"49",x"a0",x"a0",x"60",x"80",x"40",x"60",x"60",x"40",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"80",x"80",x"60",x"60",x"40",x"80",x"60",x"60",x"80",x"60",x"40",x"60",x"80",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"40",x"60",x"60",x"40",x"80",x"40",x"60",x"40",x"80",x"40",x"60",x"40",x"80",x"60",x"40",x"60",x"80",x"60",x"80",x"40",x"25",
x"49",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",
x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
x"a0",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"80",x"a0",x"60",x"a0",x"80",x"a0",x"40",x"49",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"80",x"80",x"a0",x"80",x"a0",x"80",x"60",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",
x"80",x"a0",x"80",x"a0",x"60",x"80",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"80",x"60",x"a0",x"80",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"49",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",
x"60",x"a0",x"a0",x"80",x"80",x"60",x"a0",x"60",x"80",x"80",x"80",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"a0",x"80",x"60",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"a0",x"60",
x"a0",x"80",x"80",x"a0",x"80",x"60",x"60",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"60",x"a0",x"60",x"80",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"80",x"40",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",
x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"60",x"80",x"a0",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"80",x"40",x"80",x"60",x"60",x"a0",x"80",x"60",x"40",x"60",x"a0",x"60",x"80",x"40",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"24",x"49",x"49",x"a0",x"60",x"a0",x"a0",x"40",x"a0",x"60",x"80",
x"60",x"a0",x"60",x"60",x"40",x"60",x"60",x"80",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"80",x"60",x"80",x"80",x"40",x"80",x"60",x"60",x"80",x"40",x"60",x"80",x"60",x"80",x"60",x"40",x"24",x"49",x"49",x"a0",x"a0",x"60",x"60",x"40",x"60",x"80",x"60",
x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"49",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"24",x"49",x"49",x"a0",x"60",x"40",x"60",x"40",x"40",x"60",x"40",
x"25",x"25",x"25",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
x"49",x"c0",x"80",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"c0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"a0",x"80",x"80",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"40",x"25",
x"49",x"c0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"60",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"25",x"49",x"6d",x"c0",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"40",x"25",
x"49",x"a0",x"60",x"a0",x"a0",x"60",x"80",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"80",x"a0",x"60",x"80",x"a0",x"60",x"80",x"a0",x"80",x"60",x"60",x"a0",x"60",x"40",x"25",x"49",x"6d",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"60",x"a0",x"80",x"60",x"80",x"80",x"a0",x"a0",x"60",x"a0",x"40",x"60",x"40",x"25",
x"49",x"a0",x"a0",x"80",x"a0",x"40",x"a0",x"40",x"60",x"80",x"a0",x"80",x"60",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"60",x"40",x"40",x"25",x"49",x"6d",x"c0",x"60",x"a0",x"60",x"80",x"80",x"60",x"80",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"60",x"40",x"25",
x"49",x"a0",x"60",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"40",x"60",x"60",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"a0",x"80",x"60",x"40",x"60",x"80",x"60",x"40",x"25",
x"49",x"a0",x"a0",x"60",x"60",x"60",x"60",x"40",x"60",x"40",x"60",x"60",x"80",x"60",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"60",x"80",x"60",x"80",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"40",x"a0",x"40",x"60",x"a0",x"40",x"60",x"80",x"40",x"a0",x"40",x"a0",x"40",x"a0",x"60",x"60",x"40",x"25",
x"49",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"25",
x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",
x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",
x"a0",x"60",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"80",x"60",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"40",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"a0",x"60",x"80",x"80",x"80",x"60",x"80",x"60",x"80",x"80",x"60",
x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"40",x"a0",x"40",x"80",x"80",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"49",x"49",x"6d",x"c0",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"80",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"80",x"a0",x"80",x"60",x"a0",x"60",
x"a0",x"80",x"60",x"a0",x"80",x"a0",x"80",x"60",x"80",x"60",x"40",x"49",x"49",x"49",x"c0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"40",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"60",x"a0",x"80",x"60",x"80",x"80",x"60",x"80",x"a0",x"60",x"40",x"49",x"49",x"6d",x"c0",x"60",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",
x"a0",x"80",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"40",x"49",x"49",x"49",x"c0",x"60",x"a0",x"60",x"40",x"80",x"a0",x"60",x"80",x"80",x"a0",x"80",x"a0",x"60",x"80",x"40",x"60",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"a0",x"40",x"49",x"49",x"49",x"a0",x"a0",x"60",x"a0",x"a0",x"60",x"a0",x"80",x"80",x"60",x"a0",x"60",x"a0",x"60",x"80",x"80",x"a0",x"60",x"80",x"a0",x"60",
x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"40",x"49",x"49",x"49",x"80",x"60",x"a0",x"a0",x"40",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"80",x"60",x"a0",x"80",x"60",x"80",x"60",x"80",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"40",x"a0",x"60",x"a0",x"a0",x"80",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"a0",x"a0",x"60",
x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",
x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",
x"49",x"c0",x"a0",x"80",x"80",x"a0",x"60",x"a0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"a0",x"60",x"60",x"a0",x"40",x"49",x"49",x"49",x"c0",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"40",x"a0",x"80",x"40",x"80",x"80",x"60",x"a0",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"a0",x"40",x"25",
x"49",x"c0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"80",x"80",x"60",x"a0",x"60",x"80",x"40",x"a0",x"80",x"60",x"a0",x"40",x"80",x"80",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"60",x"80",x"60",x"60",x"40",x"80",x"40",x"80",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"40",x"25",
x"49",x"c0",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"80",x"80",x"80",x"40",x"60",x"a0",x"40",x"80",x"40",x"80",x"60",x"80",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"80",x"a0",x"60",x"60",x"80",x"a0",x"60",x"40",x"a0",x"60",x"40",x"80",x"a0",x"40",x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"40",x"25",
x"49",x"c0",x"a0",x"80",x"a0",x"80",x"60",x"a0",x"80",x"60",x"80",x"a0",x"60",x"a0",x"40",x"80",x"a0",x"60",x"a0",x"40",x"80",x"a0",x"40",x"80",x"a0",x"60",x"a0",x"a0",x"a0",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"a0",x"80",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"60",x"40",x"80",x"60",x"a0",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"a0",x"80",x"a0",x"40",x"25",
x"49",x"c0",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"80",x"60",x"a0",x"40",x"24",x"49",x"49",x"c0",x"a0",x"60",x"60",x"a0",x"60",x"60",x"40",x"a0",x"40",x"a0",x"40",x"80",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"60",x"a0",x"60",x"80",x"80",x"60",x"60",x"40",x"25",
x"49",x"a0",x"a0",x"60",x"a0",x"60",x"80",x"60",x"80",x"80",x"60",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"60",x"40",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"40",x"24",x"49",x"49",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"40",x"60",x"a0",x"60",x"40",x"80",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"40",x"25",
x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",
x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"49",x"25",x"25",x"24",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",
x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"49",x"49",x"49",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",
x"60",x"a0",x"40",x"a0",x"a0",x"60",x"80",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"a0",x"a0",x"a0",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"60",x"40",x"49",x"49",x"49",x"c0",x"a0",x"60",x"80",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",
x"a0",x"60",x"60",x"a0",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"40",x"60",x"60",x"80",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"a0",x"60",x"60",x"40",x"60",x"80",x"60",x"a0",x"80",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"80",x"40",x"a0",x"60",x"a0",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"80",x"40",
x"a0",x"60",x"40",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"40",x"a0",x"80",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"60",x"60",x"a0",x"60",x"60",x"60",x"a0",x"40",x"a0",x"40",x"a0",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"40",x"80",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"60",x"60",x"a0",x"a0",x"80",x"60",x"80",x"60",x"60",x"60",x"80",
x"60",x"80",x"40",x"80",x"60",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"40",x"60",x"60",x"60",x"a0",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"40",x"60",x"a0",x"60",x"a0",x"40",x"a0",x"60",x"80",x"60",x"a0",x"60",x"80",x"60",x"60",x"a0",x"60",x"a0",x"80",x"40",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"c0",x"a0",x"60",x"40",x"a0",x"80",x"60",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",
x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"80",x"a0",x"60",x"a0",x"60",x"40",x"80",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"40",x"a0",x"a0",x"60",x"a0",x"60",x"60",x"80",x"40",x"60",x"40",x"a0",x"60",x"a0",x"60",x"60",x"60",x"60",x"80",x"60",x"40",x"80",x"60",x"60",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"80",x"a0",x"60",x"a0",x"80",x"60",x"60",x"40",x"a0",x"60",x"a0",
x"60",x"a0",x"60",x"60",x"60",x"80",x"80",x"60",x"80",x"60",x"60",x"40",x"a0",x"60",x"a0",x"60",x"80",x"40",x"25",x"49",x"49",x"c0",x"40",x"a0",x"60",x"a0",x"60",x"60",x"60",x"80",x"40",x"80",x"60",x"80",x"40",x"a0",x"60",x"60",x"a0",x"80",x"60",x"a0",x"40",x"a0",x"40",x"80",x"40",x"25",x"49",x"49",x"c0",x"60",x"a0",x"40",x"60",x"40",x"a0",x"60",x"a0",x"60",x"40",x"60",x"a0",x"40",
x"60",x"80",x"40",x"a0",x"60",x"60",x"80",x"60",x"60",x"60",x"a0",x"40",x"a0",x"60",x"60",x"80",x"60",x"40",x"25",x"49",x"49",x"a0",x"a0",x"40",x"60",x"a0",x"60",x"a0",x"40",x"80",x"60",x"a0",x"60",x"a0",x"60",x"60",x"a0",x"60",x"60",x"a0",x"60",x"80",x"60",x"80",x"60",x"80",x"40",x"25",x"49",x"49",x"a0",x"60",x"60",x"40",x"a0",x"40",x"a0",x"60",x"a0",x"60",x"a0",x"60",x"a0",x"60",
x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"25",x"49",x"49",x"a0",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"24",x"49",x"49",x"a0",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",

--Blue Stone Texture MSB = 01

x"49",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"49",x"49",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"25",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",
x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",
x"00",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",
x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"24",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",
x"00",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
x"00",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
x"00",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"00",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"00",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"00",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"02",x"02",x"00",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"03",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",
x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",
x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",
x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",
x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",
x"24",x"24",x"24",x"24",x"24",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"02",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"00",x"24",x"02",x"01",x"02",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"00",x"24",x"02",x"02",x"01",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"03",x"4b",x"03",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"03",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"01",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"02",x"02",x"02",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"01",x"01",x"02",x"01",x"02",x"01",x"01",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",x"24",x"02",x"02",x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",
x"49",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"49",x"49",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"24",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",

--Wood Texture MSB = 10

x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",
x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"48",x"24",x"44",x"48",x"48",
x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",
x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"68",x"48",x"48",x"8d",x"24",x"48",x"8d",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",
x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"48",x"48",x"68",x"48",x"8d",x"24",x"48",x"8d",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"8d",x"24",x"48",x"8d",x"68",

--Mossy Texture MSB = 11

x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"d4",x"d4",x"d4",x"d4",x"d4",x"db",x"db",x"db",x"db",x"db",x"db",x"b4",x"b4",x"b4",x"db",x"24",x"49",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"d4",x"d4",x"d4",x"6d",x"92",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"da",x"b4",x"b4",x"b4",x"b4",x"92",x"b6",x"d4",x"d4",x"da",x"b6",x"b6",x"d4",x"d4",x"92",x"24",x"49",x"92",x"b6",x"b6",x"92",x"d4",x"6d",x"d4",x"90",x"90",x"90",x"6c",x"49",x"49",x"49",x"24",x"49",x"6d",x"90",x"90",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"24",x"49",x"49",x"db",x"da",x"b4",x"b4",x"b4",x"6c",x"92",x"d4",x"d4",x"90",x"b6",x"b6",x"b6",x"90",x"b4",x"6d",x"24",x"49",x"b6",x"db",x"b6",x"92",x"6d",x"d4",x"6d",x"6c",x"90",x"6c",x"49",x"6d",x"49",x"49",x"24",x"49",x"90",x"d4",x"d8",x"90",x"6c",x"92",x"b6",x"b6",x"d4",x"d4",x"d4",x"6d",x"6d",x"d4",x"d4",x"92",x"92",x"92",x"92",
x"da",x"b6",x"b4",x"b6",x"b6",x"b6",x"92",x"92",x"24",x"49",x"49",x"db",x"da",x"90",x"90",x"90",x"6c",x"92",x"d4",x"90",x"b6",x"b6",x"92",x"92",x"92",x"90",x"49",x"24",x"49",x"92",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"6d",x"90",x"6c",x"49",x"6d",x"49",x"49",x"24",x"49",x"90",x"d8",x"b4",x"6c",x"6d",x"6d",x"b6",x"db",x"d4",x"d8",x"d8",x"49",x"6d",x"d4",x"d4",x"90",x"6d",x"da",x"da",
x"b6",x"b6",x"b4",x"b4",x"49",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"db",x"b6",x"90",x"90",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"90",x"92",x"6d",x"92",x"90",x"49",x"24",x"49",x"49",x"b6",x"d4",x"90",x"b6",x"92",x"92",x"6d",x"48",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"90",x"d8",x"6c",x"6d",x"92",x"b6",x"d8",x"d4",x"6d",x"90",x"90",x"49",x"6d",x"90",x"90",x"6c",x"49",x"92",x"92",
x"b6",x"92",x"6c",x"49",x"92",x"92",x"92",x"6d",x"24",x"49",x"49",x"db",x"da",x"90",x"6c",x"6c",x"6d",x"b6",x"92",x"92",x"92",x"90",x"92",x"92",x"6d",x"92",x"49",x"24",x"49",x"49",x"6d",x"90",x"90",x"b4",x"92",x"b6",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"90",x"90",x"6c",x"6d",x"6d",x"d4",x"d4",x"d4",x"6d",x"6c",x"90",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"b4",x"6d",
x"b6",x"b6",x"6d",x"92",x"b6",x"92",x"6d",x"49",x"24",x"49",x"49",x"db",x"da",x"92",x"6d",x"6d",x"92",x"b6",x"92",x"da",x"6d",x"90",x"92",x"b6",x"92",x"92",x"49",x"24",x"49",x"49",x"6d",x"92",x"b6",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"49",x"49",x"49",x"25",x"49",x"90",x"6c",x"6d",x"92",x"92",x"6d",x"d4",x"6d",x"6d",x"6c",x"6c",x"49",x"6d",x"6d",x"92",x"6d",x"6d",x"90",x"6d",
x"92",x"b6",x"b6",x"6d",x"6d",x"92",x"49",x"49",x"24",x"25",x"49",x"db",x"b6",x"b6",x"92",x"6d",x"92",x"d4",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"92",x"49",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"6d",x"92",x"6d",x"b6",x"b6",x"6d",x"92",x"b6",x"6d",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"6d",x"6d",
x"92",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"25",x"49",x"db",x"db",x"b6",x"6d",x"92",x"6d",x"d4",x"b4",x"6d",x"92",x"92",x"92",x"b6",x"92",x"92",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"90",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"92",
x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"db",x"db",x"92",x"6d",x"92",x"92",x"d4",x"90",x"6d",x"b6",x"92",x"b6",x"92",x"b6",x"92",x"49",x"25",x"24",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"90",x"49",x"92",x"b6",x"d8",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"6d",
x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"db",x"b6",x"92",x"6d",x"d4",x"b4",x"90",x"6d",x"92",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"6c",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"90",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"49",x"49",x"92",x"db",x"da",x"92",x"6d",x"92",x"90",x"6d",x"92",x"92",x"b6",x"6d",x"92",x"90",x"92",x"49",x"49",x"24",x"49",x"49",x"6d",x"b6",x"fc",x"fc",x"db",x"db",x"db",x"da",x"da",x"db",x"d4",x"6c",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",
x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"6d",x"b6",x"da",x"92",x"b6",x"92",x"92",x"92",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"25",x"49",x"b6",x"fc",x"d4",x"90",x"92",x"92",x"b6",x"92",x"b6",x"90",x"6d",x"48",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"da",x"b6",x"92",x"b6",x"92",x"6d",x"92",x"92",x"6d",x"92",x"b6",x"90",x"49",x"49",x"49",x"24",x"25",x"49",x"b6",x"d4",x"90",x"6d",x"b6",x"92",x"d8",x"d8",x"92",x"90",x"49",x"6c",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"b6",x"92",x"d4",x"90",x"6d",x"b6",x"92",x"b6",x"92",x"6c",x"49",x"6d",x"49",x"24",x"25",x"49",x"b6",x"d8",x"90",x"6d",x"92",x"d4",x"d8",x"6d",x"92",x"90",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"25",x"24",x"49",x"49",x"b6",x"b6",x"90",x"92",x"90",x"90",x"b6",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"d8",x"d8",x"6d",x"6d",x"b6",x"d8",x"d8",x"6d",x"92",x"6c",x"49",x"49",x"49",x"49",x"d8",x"b4",x"b4",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"da",x"d4",x"b4",x"db",x"db",x"d4",x"90",x"6d",x"6d",x"49",x"24",x"49",x"49",x"92",x"b6",x"6c",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"24",x"24",x"49",x"d8",x"6d",x"92",x"6d",x"92",x"90",x"6c",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"b4",x"b4",x"90",x"6d",x"25",x"49",x"6d",x"b6",x"d4",x"d4",x"d4",x"db",x"b4",x"b6",x"b6",x"d4",x"d4",x"d4",x"db",
x"d4",x"b4",x"90",x"b4",x"b4",x"90",x"6c",x"49",x"6d",x"49",x"24",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"92",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"49",x"6d",x"92",x"6d",x"92",x"d8",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"90",x"90",x"49",x"6d",x"24",x"49",x"92",x"d4",x"d4",x"d4",x"6d",x"d8",x"90",x"6d",x"b6",x"d4",x"90",x"90",x"6d",
x"b4",x"90",x"b6",x"b4",x"90",x"90",x"6c",x"49",x"6d",x"49",x"24",x"49",x"49",x"49",x"92",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"25",x"24",x"24",x"25",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"90",x"90",x"6d",x"49",x"24",x"49",x"92",x"d4",x"d4",x"6d",x"92",x"90",x"90",x"6d",x"92",x"d4",x"90",x"90",x"6d",
x"90",x"b6",x"92",x"b4",x"90",x"6c",x"6c",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"90",x"92",x"49",x"24",x"49",x"92",x"b6",x"6d",x"92",x"92",x"90",x"6d",x"6d",x"b6",x"d4",x"90",x"90",x"92",
x"b6",x"92",x"b6",x"b4",x"6c",x"49",x"49",x"92",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"92",x"b6",x"92",x"b6",x"49",x"24",x"49",x"92",x"b6",x"92",x"b6",x"92",x"b6",x"6d",x"b6",x"6d",x"b6",x"90",x"6c",x"6d",
x"92",x"b6",x"6d",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"6d",x"49",x"25",x"49",x"6d",x"b6",x"db",x"b6",x"b6",x"6d",x"24",x"49",x"92",x"92",x"b6",x"d8",x"92",x"92",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"92",
x"92",x"d4",x"90",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"92",x"d4",x"d4",x"b4",x"90",x"92",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"90",x"d4",x"d4",x"d4",x"b4",x"da",x"db",x"db",x"db",x"d4",x"d4",x"d4",x"d4",x"b4",x"90",x"90",x"24",x"49",x"6d",x"db",x"b6",x"db",x"b6",x"6d",x"24",x"49",x"6d",x"92",x"b6",x"92",x"92",x"b6",x"92",x"d8",x"92",x"6d",x"b6",x"92",x"b6",
x"92",x"90",x"90",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"d4",x"b4",x"b4",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"90",x"d4",x"b4",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"90",x"6d",x"90",x"90",x"90",x"90",x"6c",x"24",x"49",x"92",x"db",x"b6",x"b6",x"b6",x"d8",x"24",x"49",x"d8",x"b6",x"92",x"b6",x"92",x"d8",x"d8",x"6d",x"b6",x"92",x"92",x"b6",x"92",
x"92",x"90",x"92",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"49",x"b4",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"92",x"db",x"92",x"92",x"90",x"92",x"d4",x"b6",x"92",x"92",x"6d",x"b6",x"90",x"6d",x"90",x"6c",x"48",x"24",x"49",x"92",x"d8",x"92",x"92",x"b6",x"90",x"24",x"49",x"90",x"48",x"6d",x"6d",x"d8",x"b4",x"90",x"6c",x"48",x"6d",x"6d",x"49",x"6d",
x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b4",x"90",x"6d",x"6d",x"92",x"90",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"d8",x"b6",x"92",x"d4",x"90",x"92",x"d4",x"d4",x"b6",x"92",x"90",x"b6",x"90",x"6d",x"48",x"24",x"49",x"92",x"b4",x"6d",x"92",x"b6",x"6c",x"24",x"49",x"48",x"49",x"49",x"49",x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"b4",x"90",x"6d",x"92",x"92",x"6d",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"d4",x"b6",x"d4",x"90",x"6d",x"92",x"d4",x"90",x"92",x"b6",x"92",x"92",x"6d",x"6d",x"48",x"24",x"49",x"92",x"6d",x"92",x"b6",x"db",x"48",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",
x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"49",x"49",x"49",x"db",x"6d",x"92",x"b6",x"90",x"92",x"90",x"6c",x"6d",x"24",x"49",x"49",x"92",x"db",x"b4",x"92",x"d4",x"6c",x"6d",x"b6",x"92",x"b6",x"92",x"6d",x"b4",x"90",x"6d",x"6d",x"48",x"24",x"49",x"d8",x"db",x"b6",x"db",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",
x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"24",x"db",x"92",x"92",x"b6",x"90",x"92",x"6d",x"6d",x"6d",x"48",x"24",x"49",x"92",x"db",x"b4",x"b6",x"90",x"6c",x"6d",x"92",x"6d",x"92",x"b6",x"92",x"b4",x"90",x"6d",x"49",x"48",x"24",x"49",x"b4",x"db",x"b6",x"b6",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"6d",x"92",x"b6",x"b4",x"b4",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"24",x"db",x"b6",x"da",x"92",x"6c",x"b6",x"92",x"6d",x"6d",x"48",x"24",x"49",x"92",x"db",x"b6",x"d4",x"90",x"6c",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"b4",x"90",x"92",x"49",x"48",x"24",x"6c",x"90",x"db",x"b6",x"b6",x"b4",x"49",x"24",x"49",x"6c",x"90",x"90",x"90",x"b4",x"b4",x"90",x"90",x"49",x"49",x"49",x"49",x"49",
x"6d",x"b6",x"b4",x"b4",x"90",x"6d",x"b6",x"b6",x"b6",x"b6",x"49",x"24",x"db",x"b6",x"92",x"b6",x"6d",x"92",x"6d",x"92",x"6d",x"48",x"24",x"49",x"6d",x"92",x"d4",x"90",x"6c",x"6d",x"6d",x"b6",x"92",x"92",x"6d",x"92",x"b4",x"90",x"6d",x"49",x"48",x"24",x"49",x"90",x"db",x"db",x"b4",x"90",x"49",x"24",x"49",x"6d",x"90",x"6c",x"90",x"90",x"90",x"b4",x"b4",x"b4",x"90",x"92",x"49",x"49",
x"6d",x"b4",x"90",x"90",x"6d",x"92",x"b6",x"b4",x"b4",x"6d",x"6d",x"24",x"db",x"da",x"b6",x"92",x"b6",x"90",x"92",x"b6",x"6d",x"48",x"24",x"49",x"49",x"92",x"90",x"6c",x"6d",x"6d",x"92",x"92",x"b6",x"6d",x"92",x"6d",x"b4",x"90",x"6d",x"49",x"49",x"24",x"49",x"90",x"db",x"b6",x"b4",x"6c",x"49",x"24",x"49",x"92",x"6d",x"6d",x"90",x"90",x"90",x"90",x"6c",x"6c",x"6c",x"6d",x"49",x"49",
x"6d",x"b4",x"90",x"6d",x"6d",x"b6",x"6d",x"b4",x"90",x"6d",x"6d",x"24",x"db",x"92",x"92",x"92",x"b6",x"92",x"92",x"6d",x"6d",x"48",x"24",x"25",x"49",x"b6",x"db",x"b6",x"d4",x"d4",x"90",x"92",x"6d",x"6d",x"6d",x"6d",x"b4",x"90",x"6d",x"49",x"25",x"24",x"6c",x"92",x"da",x"b6",x"b4",x"48",x"49",x"24",x"49",x"db",x"b6",x"b6",x"90",x"6c",x"6d",x"6d",x"48",x"6d",x"6d",x"6d",x"49",x"49",
x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"92",x"b4",x"6c",x"6d",x"49",x"24",x"db",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"48",x"24",x"25",x"49",x"92",x"db",x"b6",x"d4",x"90",x"6c",x"6d",x"92",x"92",x"92",x"b6",x"90",x"90",x"6d",x"49",x"24",x"24",x"90",x"92",x"da",x"b6",x"90",x"6c",x"48",x"24",x"49",x"da",x"b6",x"92",x"90",x"6c",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"49",x"49",
x"6d",x"b6",x"b6",x"92",x"b6",x"b6",x"b4",x"90",x"6c",x"6d",x"49",x"24",x"db",x"b6",x"6d",x"92",x"d4",x"b4",x"6d",x"92",x"6d",x"48",x"24",x"24",x"49",x"6d",x"da",x"b6",x"90",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"b4",x"90",x"6d",x"6d",x"49",x"24",x"24",x"49",x"92",x"da",x"92",x"6c",x"48",x"48",x"24",x"49",x"b6",x"b6",x"b6",x"90",x"6c",x"6d",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",
x"6d",x"db",x"92",x"b6",x"92",x"92",x"90",x"6c",x"6c",x"6d",x"49",x"24",x"b6",x"db",x"92",x"92",x"b4",x"90",x"92",x"b6",x"6d",x"48",x"48",x"24",x"49",x"49",x"b6",x"db",x"6c",x"6d",x"6d",x"92",x"b6",x"92",x"90",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"49",x"49",x"6d",x"b6",x"6d",x"6c",x"48",x"48",x"49",x"49",x"b6",x"b6",x"92",x"90",x"90",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"49",x"49",
x"6d",x"db",x"b6",x"b6",x"92",x"92",x"6c",x"6c",x"6d",x"6d",x"49",x"24",x"b6",x"db",x"6d",x"b6",x"92",x"92",x"92",x"92",x"6d",x"48",x"48",x"24",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"6d",x"db",x"b6",x"92",x"b4",x"90",x"92",x"6d",x"92",x"92",x"49",x"24",x"92",x"db",x"b6",x"6d",x"b6",x"b6",x"6d",x"92",x"6d",x"49",x"48",x"24",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"48",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",
x"6d",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b4",x"90",x"6d",x"49",x"24",x"6d",x"db",x"92",x"92",x"b6",x"92",x"6d",x"92",x"6d",x"49",x"48",x"24",x"25",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"6d",x"db",x"b4",x"b4",x"92",x"92",x"b4",x"90",x"90",x"6d",x"49",x"24",x"49",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"49",x"48",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"90",x"90",x"90",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",
x"6d",x"b4",x"b4",x"90",x"b6",x"92",x"90",x"6c",x"6c",x"6d",x"49",x"24",x"49",x"db",x"92",x"92",x"90",x"6d",x"92",x"6d",x"6d",x"49",x"48",x"24",x"25",x"49",x"6d",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"d4",x"d4",x"b4",x"90",x"b6",x"b6",x"d8",x"b4",x"b6",x"d4",x"b4",x"90",x"b6",x"6d",x"49",x"49",
x"6d",x"b4",x"90",x"6d",x"92",x"92",x"92",x"6c",x"6c",x"6d",x"24",x"25",x"49",x"db",x"b6",x"92",x"90",x"6d",x"b6",x"92",x"6d",x"49",x"48",x"24",x"24",x"49",x"6c",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"90",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"b4",x"90",x"90",x"90",x"b6",x"b6",x"d8",x"b4",x"b6",x"b6",x"b4",x"b4",x"b4",x"90",x"6d",x"25",x"49",
x"6d",x"b4",x"90",x"6d",x"b6",x"92",x"92",x"92",x"92",x"49",x"24",x"25",x"49",x"db",x"92",x"b6",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"48",x"24",x"24",x"49",x"6c",x"d4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"b6",x"b6",x"b6",x"b6",x"b6",x"d4",x"90",x"92",x"b6",x"92",x"b4",x"90",x"b6",x"92",x"d4",x"d4",x"b4",x"6d",x"92",x"b6",x"b4",x"90",x"b4",x"90",x"6d",x"49",x"25",x"49",
x"6d",x"b4",x"90",x"92",x"92",x"b6",x"92",x"b6",x"92",x"49",x"24",x"49",x"49",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"6d",x"49",x"48",x"24",x"24",x"49",x"25",x"b4",x"b4",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"6c",x"92",x"b6",x"b6",x"b6",x"90",x"90",x"b6",x"b6",x"92",x"b6",x"92",x"b6",x"d4",x"b4",x"b4",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"b4",x"6d",x"6d",x"49",x"25",x"49",
x"49",x"90",x"6d",x"92",x"b6",x"92",x"b6",x"92",x"6d",x"49",x"24",x"49",x"49",x"da",x"92",x"92",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"92",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"6c",x"6c",x"6d",x"b6",x"b6",x"b6",x"92",x"6d",x"92",x"b6",x"92",x"92",x"b6",x"d4",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"92",x"92",x"b4",x"6d",x"6d",x"49",x"25",x"49",
x"49",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"25",x"49",x"49",x"b6",x"b6",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"b6",x"90",x"6c",x"6c",x"6c",x"6c",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"92",x"92",x"d4",x"d4",x"92",x"92",x"6d",x"6d",x"92",x"92",x"d8",x"b4",x"b6",x"b6",x"92",x"b4",x"6d",x"6d",x"49",x"25",x"49",
x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"92",x"92",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"da",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"90",x"b6",x"b6",x"b6",x"92",x"b6",x"d4",x"b6",x"92",x"92",x"b6",x"92",x"92",x"92",x"b6",x"b4",x"90",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"49",
x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"49",x"25",x"b6",x"db",x"da",x"6d",x"6d",x"92",x"92",x"b4",x"b4",x"90",x"b6",x"92",x"92",x"b6",x"92",x"b6",x"b6",x"b6",x"92",x"b4",x"b6",x"b4",x"b6",x"92",x"b6",x"b4",x"90",x"92",x"b6",x"b6",x"92",x"b4",x"b4",x"6d",x"49",x"24",x"49",
x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"25",x"92",x"da",x"b6",x"92",x"b6",x"92",x"b6",x"b4",x"b4",x"6c",x"92",x"b6",x"92",x"b6",x"92",x"92",x"92",x"d8",x"b4",x"6c",x"92",x"b6",x"b6",x"92",x"b6",x"92",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"6d",x"49",x"24",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"90",x"6c",x"6c",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"d8",x"b4",x"6c",x"b6",x"92",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"92",x"92",x"d4",x"92",x"92",x"92",x"6d",x"49",x"24",x"49",
x"49",x"6d",x"b6",x"d4",x"d4",x"d4",x"90",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"6d",x"6d",x"6d",x"92",x"b4",x"b6",x"6c",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"49",
x"49",x"b6",x"d4",x"d8",x"d4",x"d4",x"d4",x"d4",x"b4",x"90",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",
x"49",x"b6",x"d4",x"d8",x"b4",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b4",x"d8",x"d8",x"d4",x"d4",x"d4",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",
x"49",x"b6",x"b6",x"92",x"b4",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"49",x"49",
x"49",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"90",x"90",x"90",x"92",x"92",x"b6",x"db",x"d8",x"d8",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"d8",x"b4",x"90",x"b6",x"b6",x"da",x"b6",x"da",x"b6",x"b6",x"d4",x"90",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"92",x"d8",x"90",x"92",x"6d",x"6d",x"24",x"49",x"49",x"49",x"90",x"b4",x"b4",x"b4",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6c",x"b4",x"90",x"90",x"6c",x"6c",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"b4",x"90",x"48",x"b6",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"da",x"b6",x"b6",x"b6",x"b6",x"b6",x"da",x"b6",x"6d",x"b6",x"da",x"b6",x"92",x"92",x"6d",x"49",x"24",x"49",x"49",x"49",x"b4",x"90",x"90",x"90",x"6d",x"db",x"db",x"b6",x"49",x"49",x"90",x"d4",x"d4",x"d4",x"90",x"6d",x"d4",x"b6",x"b6",x"da",x"d4",x"b6",x"92",x"6d",x"49",x"49",x"49",
x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"90",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"90",x"90",x"6c",x"6d",x"b6",x"b6",x"b6",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"92",x"d4",x"90",x"6d",x"b6",x"db",x"92",x"24",x"49",
x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"b6",x"90",x"6c",x"6d",x"92",x"6d",x"92",x"92",x"6d",x"49",x"92",x"92",x"b6",x"92",x"b6",x"d4",x"d4",x"b6",x"b6",x"90",x"90",x"6d",x"92",x"b6",x"49",x"24",x"49",
x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"48",x"48",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"b6",x"d4",x"d4",x"90",x"6d",x"b6",x"90",x"6d",x"6d",x"92",x"92",x"49",x"24",x"49",
x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"49",x"49",x"48",x"48",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6c",x"48",x"49",x"49",x"49",x"6c",x"48",x"49",x"49",x"49",x"49",x"49",x"24",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"



);

begin

process(addr)
begin
	
	data <= ROM(to_integer(addr));

end process;
end rtl;