��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ��>�(Ŗ�XV���=�<4����>c���t����֪� ��?��A������.�.��G� ��{~�޻9zZ��/a���<A�Q%�W��F�8�"�uRȸX*�V@��L���uZ�5t.yѤ���lN�t(�����.�}��
�9r��w�R��}����\qDu��d?e��r��y�ޣ�y�$�5Kȕ�7O�Q�g�������R�ɧو*B���UR<��5;_n���ݵ9,�!��*�w����#��t�0ߠDS���g�.Q#�S���b#it�`B{3�����)o��Ǉ>��~���ƉK���4�1Vq�"Ӹ��7ŤN
|4��7c�FM����f��=���#ݡ�<\��N볕Y���Uo����Ol�~�� =z��S��mz)79�v�t����K�p){o��%���ʚsj}���ʾ 4�)�f��+�:�H�]�$~;W��[f	4|�������o�h���{58�FmpXr�8�	�����D}CNs�{Ε��7^"�ن"�/��	�$'��\3L��d}{̻}�����kM;�h��C1�lV��cq�w�/�
���$�����(o���4}��nf�u+��'�/��|gK�I�l��6wY<�KjY\v�gզ=f֍��"]�_#Lr+p��b�ȿL7Sp�"H#�M�������da��`U"����070��\�*�b@������dd	��c�sv"t�!�sg_N�e73T��t����m���E�-�g�&����\=D�8G�uвyQ�}�����i#�x('��{�sO���;@m��֌�G�Ka_��.sWʵ����b��v��(�MzP0��t[t��f��I�%��� ����ֺ�e��^i�"v�n#��Ʉ%}�_�IY�B�7�,ǖ�^d���\\у�^�Rl���9�1P2Wa�e�ޖ��W4�Lj� ���B�쏄׷�2����]����؛�h�\�8�������e���܌�8��ih�i��1�JF�mɍ�z��� �Ӯ��;1�n�E��<�:�=��y���7��]���]��V���J#\�p8�u4�>w��Դ����#�I���EA
�5�q��8fmޞ�����ʜ�6������[���!Tc
:*<힚���K���=yEvg���6�(��3]�ޅ�>P��p���ߐ"��E.�5Ar�0ᥘFj�v�}��+1鬌���h�n�.kH�!��<�nk.1w�_4�'�i	��CXN�s?��d�����.Z��`�厗ܧXHN�	��{��bZ�9�L�4��xbx�ݳ
i8[�u�y���V��Xs�hc�q�O��F���o�!�uM��8֫�ƥ>A����0<���8
 ��ab�xz�.0M����Zс죄��*�����D9�:����;�\_d�<u�y���NUBD�JAna|w>��d�A����oK���v��јp�	ۢ�x�Z�����KHU.�Kȉ�>q)���LQ���Srx�׺:���P��^�	I���{��z/E*UE��K%���^����GC̒#16�D��v��	cY��J�p*����#z0�>u96�0]v��ipO�s�K�Ql����c��>�E�H;g�{r���h'��h�`����Qf6T�����Ho��,���D��i�R�B��ՀH�e���	�飓��4y>��+�U�����.���f�z:�����a�&����>���ڛ�/���(��yX�S�/P`�ՌK��F~[�ᡣ����.��(T�S��XujB�������(=�}�%x+��k����:��phA?hVv�
âd)�k�`%ڳ1u�� ���Gd�,��6���%�|�QG��M��;�P?�#�@����(��K�|�0Xz9��H�m!��iM�W�����$t�K
��.�>�L�gV,C��.B:s������n�j)�.yO#�,�).��͓�gD�Q�ׇ��6e�c%��h ��/�N1�O�к̆��p�櫳��dR=/�����FR�L���S]HTIH�m��6�N�r?�׹BWR��
��ا�ɭ�3Z���\8"^�il�a��*���G�{�HI����
_�ސ3��<a⣒eaYS�p��#��� �ٰ��{�J߼A�(AR�-����K.�����vUh)d1y"yM3R�/�����|v������;�mU`R��U�\R r�b��J|��yGе)Kй�S�W:�ɕۛ#��އL��⤝��,�+�=R����i��R�H�p�ѽ#�BqE< ��!	��5-7��n�ݏc�1�Nx�Mں�,�� ��<dhg6�1)�g�̓P���+�^ԩZ���À'���S�������`9K��:���'��[&�rѥD�z6�@n����ܲ�I4��<�ϗ����A��n�q:g{y�����T�B�e�1>h�X�k������a�@�5�����#),�F�N ��?�C�c�aH�'��$�>��KU�+���������&�ۯ�����Nڜ'1o+X�c|�BO@�g����鯈M�%����t�X��(5����=7EC�>�Z���ʻ��B�^s�JMbF�G���l[�����T�D��2�ih��s�t�ych�� ��rGaP�R����$�"S1X7���bt���U��c8l��I��s�O���팙�]�Z����=���3A�,G�W�K����关mG[�ZT�-�&)<���E���4/����g{�7o�k�T�ÊS0�'�g��Lyu����ze�9��3gn�;�B0���2'�a�C��5�|�/��}�@�������Ga�G'=Νm.�?���q�
s�|t�}��Za�,���Ee����5�Q���b|m���u�8'���2MQ�jw롐�8G�8�^�Э�0��4�Ȩ-v�r���v�	�K(�{�,P�I����+~�74^�0
��wb
]	�j�����O<u~t��� �0Ϯ�$�����U�cƳ��^���6q2��`��hZ��	�h�����b�ٓ"��6E`xlq�u6��:Y2��m������j�E\���3���2B(�C��\ǧ����~}�����S�+��C��$����k��.��k2s���A��J�U.}(��ᆃ��fPd��E�;�D�w��l�՟6�-l���ls�4?$��Z���7o�w���r�p����X�8�qc��<��oAK�Т�^x��[z���	l`���Oző��{�RJ��(5`G?&���X9~��,r?�	�����-����g�@�+�����y[�-̹J#~���}p�Z�O�.4i�����O�-�wf��;�2�h�^�c�߹_����y-���υ����T�Dyɮ)/��A�z.�g��h�k�~4~Yصw���,�H,'*�ծ�ƙ��D3��4H(0��'@�~������r.V]#�c}P�����lb̃x�JAM���QhKJ}�����F|�i�j�<P8�2(;@�����4$u�����[h/ �墫2ί^�5Sƭdt��g|�i��0��"��p�6.����������TDj`@<���xV��d6������j�3c��j��"p���4T/J�
 ��U�Yf@Q<*O��*��΍U��<PE�Ø�:�!|'�ʔQ��� ������q���4���LMЪ�톖^4yۉ��y�?���6��D">�A��71lg;&I�(�̴��a���W(&)�� �ۨ+1)9�6��'�+����V�剙.�yf7Z�dl1N&	�t��!��L/8\|�]m��j�TR���&
���6%�1��nò_�a��$F0�8�x�0K��Z����a�-Z1����>\��w�9.���ɽtq�c�����,n%�Y�hvQ���JX�����c���M��6�.��0EM���*,��$cE��_m�8suxV �~J|�<�{-�8~
%q����;́�N�{7��e+<ÿB0-Z�mֳ���ʐRэ�<�v˔g)6{ 3R�
!�Ί^���#�©TfͰZRn�5f�	@���~͉�,��7-�[�-j�^�E���]���L�pȗ�p�)����-�e3eT�=U��S�����"dxWDj2��F�YB��S�IU���J-HˣxX�3���BJ�C;I�^�3T&N[W��̳j<c�l��!��,7��=2��}7ڥ�X�[7���SK��T0����r)��	�_@�Q`Y���K|��f�y<[%�wqz���>mYF�xg�����ʄR��p�)�"�#8��%�wM�N�g�!������7���n��խ�g\a�׆����U:�>�����~Jg�f��9��7W�g�^��|Z�Gj����ظw�툼{2I��*�;�H�9��3[�4q)W�K�]�^�p���nD�}��Nj��� �	�ջ���2��Kz�����y�9���;{����g^D��[�Wu$4�/�!7��P�A�saG���ϗ:$�F[�5�F�T��!.=�&s�o������ղ��t�nv�q��.,u��S(++i�������l�1:�|o�٫J���6�q�՚E����?9��Lw@t�I�LYն�y:ܡ�+���s��Z@� `��^��7�4P��n�G@�^�e�tXU�
]��ǜOB\^P~8u��V���ꮄ�9�T�e�����z.*����6D]��7������Zw��~�n� �4�tm�0��uٿ>��&�)O�0�)Q���5�/Q:�K{�4�R^����Jz!B��,F0��G=��8��c>Bb�\���`��	G������V�߮/��,S�\D����h�]B�(q���u���9�Q&� G9|[~��j�q:5yD�)a�0��gu�0R�7��ﳺ���A�-Gϱ	L���ag�s�ʴ�j&qpsd8q�~u&�H��̞�l��Ԕ����h���i�g�F��`[�5%t&�T���P%����.R�HI%Ǌ��<>�1ٔI~�[Y?Pb^�h�TF��3C��i�|%���[��ٹ�Q�qp������@M((�Hn���g�G�:b 5���jOg���x&g-�s׹ϛ��:�#v8嗉�;��bNr>��r���e�9{��8roS�nj&,�1u���uJ���'���P�5�e��paG��0��d�m{ܖC��ݕ���uV,g�<�/r;.os+'2fi`�}��7ZN�rG�a�yB������5/@�Vi�;�D���2��)� >
�%�.�eٛ�jߕ��D�=vO���w@X<wL������y��5w�,q�^�T�F�C������x�򉮹�_0�I����հ(ݴۃgc��L���W>���K#�����I$˛��ٵL��{��rs\������9� #�;�1���B���H�j��+]�	�CQv�N�4Kh[A���4�ܟ�w�:��2�oq]�=��oihI�ܻ�2��PvR6*:�s;orH.��dg���y��EA"�"����p�(��{��$PƉ�g����f��4���3�-�ۛ��[l)������EV3�Oè)$VB���r��}m��m's�K=>
�����+�3:�" ?	p�<�ZWD�������qlc�PYRI�\V�-�p��
��[2��q
��o%��Pi�.��_�&P�w��p�= �ہ8�+�K�{>��9�z͙�P��nƦؘ׆/������}�k��ad�n�[c� s
(�% W�C�Lg�[S_�>�]�
�{MFxr���I(�r��J�q>c����x�0�p=\�c��I)4_���t�t¡W�r��+��h�\�@H-��I�Q.��ضx�&��A���t�^	p��K ��[�������X�}sn�L�*�u�X&��7:D/f�����{�͟/ݎ�4^v &��Ix�6�����ǅ̦"�d�0!}��Lkf2�j��=4�x�7k?�)1��ぁ�=��?�;� ,=�%j�쎃��ǀ�����m�h%wX���[\}ٌ:y3�����o��u�!�O�y ���3{?�1�1aݝ0��Ff':����`ӗO�>���w�����)=�}˸�6Z~�9���Uj���VR�t�P��1�	�)��k�;�OU�,�}�S���&U�Q�#?-��^��/E�g(,2g��0���|�o�/�>����!�B�OPD�h*��tHCD����8�^�N>at5�F��"A���Vڭ����o����U(���u�F����׹v��s�/�
��Y�)��Yʑ��xƒD��q���g�z������3Q���P�q
j$=sKT�M<vp�J6�A��(�l�g�ɝ����+��2�{��@h��]�i��1t�>[?���ם9K
$w���|��[K�?��%�+��IIr�;��s;Z�ke�T5W�)��+����"V�I�����b�NTqq���+X�J�z���P[!�X��J�Ffi,&���X�/)s_����f#=F���@�f�N9����>�>	�-�?Ud�4���3����>B����%�N�W� !f����l��OcY��8M����m̥��3��	���5O�Y�f9əP�����x��/�P>6�,�s�
)�#n�Z|�3fN�!netؔ�F��["�8�K+��ٞYy=���2y���:+�r��2}�3�`{��|��	!J�*��-6ݕ��m�k��	0S�l;���ʲֈ1��7v�[��Ew�S�o��UåS{Z.�>L�$y�d���5g��H��:M�HK����:���/���K�
PJ��U�I�F���B?��Y	ԭ��d���e�}�ݨ��M/2i~7�_U��׽'l����kE����(���]���3�.Q����j�E���䶜b�팧���K��|`fYY�"�D&��9��{��l�_������%��^�a}x%F�},�:�;�ӛ3���M68�j� ƫ͌8\Gmha\Qt2�1ʷBY����9V6-�*7���
%�S͟]��b��)�uX��2�Miz�a
$�b�`8�S����`RQAp'���dS�!��/�ʤ& E����'�lin5���2�x��G|nцjP�i�|�(�HM�qh]����;�6˷᥮G��_N�/�|)IS�~ߩLR9$�KK�qZ7"|!��#H����-:R�{�� ���A�q��R A+⢢�$��M��8@�F~����v55�JG����N�>�r�ݣF��L��∬KU!��
��6��
˦��(9�Rl-���D�j �5��s�E�<��`����c����;��O|�|��Ĵ�a����i%�?{��㉊�as I29�:Hj #|���F��11����md�Kp�Qσs����\S~I�P�w���j�S;�e�7Fa4(�<�ƧRWN?LP��q�W�N?���ُ����.�O���nS��6�.�"���K���o�$D�cҌy��
s�r�@����챜BbN�^~�(=³��	��K�w7��豦�����}z�����"�	-���@�;\h=�
�n#��x�2싘�?JC|��)&<#��a�)����[�҂���  0�*�3?=��S��t�U
q$�R��V{���r�(~0D�!�@�BS~Ȍ�����&=�x���l�vwk�Jj{p�S��"	�����>����1�L��湇�`���֢��9t�Jp
�D�/��~�8�9���h~Eh7������sӾJx��ȣ*[���ԡK7H����0QE����ןSkF�w^�Bc�y��3<��[�&�Q�g�o�N��ׄ����t�iެ��M1S�]]F�7�߲UM�k_�q�$������(�Qދ�0��>�e�2�Q��7�vDh���`<,Y�hd�y�F�����|���F��Z,�B��q+6߄�R%��Ǝ�	�������*��cyA_Ti�jP$�W�b|aKô��ᾭ��0��Z��f�֠P;������ơez��V�&m�ʤ��S\�K�?É�1P�k���05�H��A�d�a�O������K8>'׳޴�.���b]��W~�Q�\�a��� <�TbK�P��x 0���ﴳ��&cQ/1o��w�j�7�u�x�gL�i>:G}jr��T�T(1л�Ld��#�a��n���Y�1&eM�Ę��,��m&���`6%��'��]qF �G�ڰ��tE��$g`yі�C��0���S{�3pX$(��n��XiIؿ	����-�(�4$��O:���$���MLҿ�B���׽Y����@�����(�U��`��{��Q�Y�T�ř,����M�Ϟ���clʗTXU8���w���	�o'w���10�tU<q�b���=�^���s�h�O�Ĕ�M.�&��XtS�͍U)�L�X/M�	�ە'A`�o�O�d�u!�R˶].sO���f$=OV}� ��b�q*��gÄ� ~�E=BW3p��}��F&��˄�>����72��۠:L{�龎�y��uq�4Gg5Cs��F<�ט�OѶ�#Ƌ�����������	#�g��ƴ�����JF���!��z�Ι����Y�-wdAbU�q�Wv����X�W�?�!�R
J4^&��aq��³���%{$H2f��	u�l���;���G�h�U��-��YEY�r���ĩ?�s�J�y!���)�#8X7�s͆�j����F)�j�~8/8k�t���9���­��l�Q���֦���I�%/�u=�R�l��[+@���1��S�s��
�5�W9���h�t�>�=��K��t��� �D#62��� ����#eVƞ*Er��a����oV��n��g�'\��UPW��N�zo�mf��\�	��H
҇��F����U���x�O�)]O��7�%Z��wgNB��'�o�I�� ���z�����^ü���^F�:�3�",���+<��t 6�S,Z�EZ��h1A������`82�wZO����>���M�����v�]|,��
�Q�����ߓH(��S���BbQAf���~d�|0�p�u��\��&���J�xH�I�W����<[5I�����5�r)��h9>`�d;���-�d_��U�����]v;)�����ǫK�f����G�*.��O�[;�O���-s�4G��J��z�ݳ�D��}���Ӄ"�DĠI��!��h��z<�~�B���9�xѐt4qc3>@%R�=-K�'>�@i��_PM�";紁�J���
���e�*q8+�{�Z�)���G��%���R<G�ivw� ����d��?�p�_x���D�ET�m���ڧd��G��R�]����#7y&���,��B���_o*a��^�~q0c���z�ة�s`��bK�J��V���-��������ߝ4���ѕ���M�aO-Y��KE��J5\�0-GӜ���긕_�)�@�9K*�4�*������y`��c/K:�Ix-�+t�rt,n��䌟B�>_7��k2��Y������\�d 9}L�o��B�)��/^�xE���&�!v� �h��JW(F��Ajԁݩ�X�8|uk�Tp@]��L��V_��[HUuyL�`)rt�Q����5�S�Q��?X�0F�Ʒ'��?&�6.��d3�#��M��p��OZ��~��)�dDwz%T����YB��z܈\��@�n���eخ��A˫O#?zlޭQlO�Q4~m17�BM�7�i"�w��������;S�e�R����S����ޞ`%?��}�o+�fӂ�pS̯��{2>����z�Z��4��bLˮ�ؒc�0+��lS� 8���t��
�����|r�UL_�+��?�{~С楱~�|SB���˖U���bց{rֈ!�ZmK�`Z9I���rP�!2�Z��ma��B�y��z"8���2�;&�N658��*��@�������&�(�B��O��p�wʪ����
��\8�Q#h��.�q�C��j���]����l������;K	2[6��$D$QH��il��`I�4�v���:�-K	\�`�����*���j����7>������8�u���o���t���^�g7�*.����6V����pSRd�X&��2m#�M�Х8�p#���̹�4��Y�J�C�e���;&
\�Y�Lۄ(�m*��?) o�R���S\��p��|�"8��3K�f���WT���YB��F���w��'�C��,��#g�����`2�h�[�^2�r���I��s4V��?��#�s/�U��7�{��1f��S1o�C�*Yk�$�����Ҋ}iԶ����+���'��U3�t���Û���y2gj����[� ��)�N��[?�2g�����S��@��RF׍�v���oQ�t3(�S�U���mX~�����Q@�׻��qꚋ��t*p�r�$}|h_)�;�L'̀�����_���D����Z���>3���lD�r�"R�/fg/ZFt��W_�����3�+�'�U�Kv1_��&�/��76r�w�wOIA�Ʉy�������}K�F�҃y�ɴ~��(��R��/�,v�"��u�Z]�L�q3�8Py�I,Y_����S��}��e���8�4�;���h�p<�"N���YgMF�bZJD�~�đ��4��pRdӴAH.�+��lϨ)M"^�j����q��`OXGu{?ye[>���t5H]�V؃�"��̍?�����&�ԕ1��C�'��^ډ?`����KEњd^f���VAΚvڪ}��0��Xf�^����&������bU,���|�t�����N���W};�e8o3�i���=oE�.�[	�e���G����w��T$$5����\�	9���n�[���ԇ(ru�Y��Cp(�
z9���|�X�]L4�*Z� !����~Ԛ��ine��<CV�vsk6D�֘z:g���b�3ϐ��ȟ��Vd��
F����Lv�r�n����P��+D���k��s�ȣ�sF�����6�OW���$ �|�'̆��^HS?+񣰍Q����r���N�Ο�׌`�y8���VAēD� �i��,=)����L����lU�E��@OF��~�Q�fd�Q!��P��J��>3���;Ϥ����(��"�@�u����,;�*�E��A���&T�Cq/5)̽mLU�{�9ڠ�ޗ,��KS£���ŀ���e��I�:�9�� ́ �4�O�Gm��!�r����nC�'#A�E�]&	��w����~��r�#��@	Q�4Ǧ^�ϻ��چ��I�@����l��?l�N&�݈:���ƅ|����������3	+���Ҧ�H�..��"z�ZHZ����	n�����+?ր"+���_l������v{�vQ�����Ox���HE1���,���hm�/4x6��w��r�Ro��EU������W9>��Qe������̵�M��X�ء/��&�gsI��>Ȏ^`�>�9�%�̦�!!d!^���x�T�Q�Z'�r��XX�8��C�V�ߍ<��8���h�X��E%]W9y���D���������rz(�Ϛ�0��l��7^dD1&[K���F���Ƹ�0��.M�=ķW�b��f��L��PY�b��Wُ��O�g�0����u�8�YD�&��j� 7�{0=f���e�p�W�j������>�g;� ��u]���h�'�+~�b�$������n��w�1\1�5t��ǙgѬ���BV�=�?o� ���3�a?�HmB�b�(-�Zgvت��=ͺ��Vw�G�`w�0��t��LF6�?�}��@��?�<�l�F��g�*��� (ln����n:��u&c/F���.����%��rB��{<�sگ����/�k�U�3Ӫ9��|�۰�T:�#��~���ש�{/)�¡h
�x�F�︟3���`(�q��bu���Eu�*b��t�rb� %"Ra��O����r������4�NГ�7m�i�f#�`�]����`P��y�� �[�����x���֛�'Pj�+���F��K�.�ѯ�����)�;��4��8#��Xg/���������P�&��q䕦u?r��)�����d�*g�g������rrYB���������q��-����'�W�*�{��U��z.�pks��ɱ��X�,�u��Ȩ���ۋ;	ћ�Yߖ�!�\��^y=���a�2�������-�kЃ��ѕrD�0Ѵ�ch�n%�B�y7R�E�x?�<2O��<,E0q�!fȺ�k�A=�H�U�1�$��||M���? :J񁅶0RO:X$�j!]8��T��q��|�(i�^~����;D*��zQl�u,	Z��\C8��Nrc�~�Gl� ���̆���?J[Ae���D�k:��rg�����6y�jc^bѢ����5���>�������{�E�
�������������=�5��H]��)�2%��e�׋�=���!�1 ��$p}�HDp��ꥆ�Y��)Wp�����W��_�l*'N�G�_m�qC����p�����J91 ���&��a�ˣ�;` ]��M�H�����}����}��,��d����S���oј.ˍ�f��f���?l;L��<����߼��W��������7\��1
�;�H�\�ok���Y�����o��$ ;46��'����d
[���G��w�`5D�ӵ@/�NM��r,�X ��^�
�#]���^���ZYt}Tt��A ��Ih�v�Ƙ>�Z0Q�חa�,�1�Z5n�[�@�.���݄��hu7�@c�4���N_��1�3��&�]� �3�c4u� ��ONVeY��1�\����N�Y��p�����C}�L͵_��x�rP�(�7;iO�e: ��10LCNVD	��!��F/Z��rP������LFZ2�4�{�u3�m	&�׌N���/�C�6#!�D���'v?*����5�}h�u}�n�oM��O<�u")�j���WQ��1#*�W��!T�����͡AB+y�:�"��IW����>�v$���?�G��Fh�Q3��������=��\��b��60L:���}@Ȳ�G70!�t
����FK�SC�RQ~��P`�k���wn�}�JG�/��J?S�Mj�+s����'Lv�'����v|ۓx��N�R2�êC��{ x�dO����������P6*/!o����wQщB�!<ɛ���gЋe�2�ۗ���J��	@l�x�������|է�R�+ʥ��?�x�S��8��V��}l�"�2��( l� �w{Z�Xݐ-yT��Ĺ��r3&�^��@M1�Z��ڪ�~�-P�-Ft���$�J;���� <1Ŋ��H�ˤ��%�CZjs9rr۳���B���@@dE�R?S��;s�&�˺�v̚�>,ߥJK�����>M�y�z�_�o�����}��ťe��y�Uz��G�\{o��	c�<�DOqi���wIB�F���iq��S�J�8Y.$!^�1��^3#7�$���?|T����gu�"���c�f��)v}�E�n�O.m��Z5$��PT"L]D�]04qn*"�j;��I�0���q��#��N)?!�rs�ګ�O���]3Ky�OW=�8}�����w3��YR8�ڔ{|k�0��;%j<N;�I�CV�P��RPC=c)�w�>A�`ǐܕ���O$�=� �|���5j�8A 1=P��ƏT���T|z��`�	g�(�6`�9��As����a����f�S�N��p�ɝ(xFK��㧾��4۬ե�F	Q�s\������\0&���|��3U��8t<6V�gKƕ-r%Js0�g�{ܑC�P����$O�T(�<W~ˍ%D�������T�А��k�M�RX�h�;*څd11\���i|Z������LRĞ��k����O�<gސ��PH�+�.VE���ń�S������G���E�MFہ,q/�D�b�&��)����z`;�����5`CJf���J�iE��eXn"����FŘ3�b�xZ��c�(��;J��h�����,�z������J4��e�3�$:ӯH� Y=W��}x��T��)�@�O��(6��&{���u#y-1�fٻ�ܑ�b�"E�W�`�
�������ӄl�L���[�Z��{�{PP�JZ�\O�z���OP=�����z��GXf7�TI����r,Z��V�M�����G�'x�l�q|��1�K�����M�_��k��.�y�P�>ɉ��OG,َ��C�$O��:X�et�Q=�΋�)�����n~C���2K�jz_?��`�6A�=�h}z�$\�#f>����F`�Ϋ��2�CKfՈ��l]�s�9Ņ�~�F,�$Z"�_�� �����bwk���j�iǠ0��:nN���Cb�gp�W6�� �	T��s��=�l��F����m�O���.�%���3ȝEQe���!:�p��Fy�X�Z��W��\��q�c�,7��l��}Fs��v�X5�kxA�~�.oCyB�}!N��r�����������(6�B��d���q�*�	�!��+Er��3�?@�Õ	�̄��v0M��Y��Uw'����~+�;8�@���3�0"�k��f�4�89�xǠ�wW��𧇽;A*��t��xx���n�"c�p�K����$��������
�X�l�w� ���H*�?��x	��Ձan��l�L� ����9�*7"c$sު;%����G�ɍ��<�y�(�?%sc�l��Fg�\���;p;5��D/���S����d��X�S�H
/s�}�|L��#�Fa�FC�LO�sۛ�����&�¸]�g��� ��|7�0}uF�ۚ���g���M���TR��b+F�����c�5��D>�<Y%����,��*�h��f����k4��R�p7F��3�ټfhz�_���_���/����
���t������,�x��\�S��܁\��z�?��r�Q��t���������l�R(4��V�(�ڵ��tA�엘��8G2%��F/�~,=\�{�gD>f۠`�5%��<�x��d�tl�z�=��ݩ��՟���,��Mr��鎠�^���1�),�F�&��M�Q^����
�r̯+��K֗�X��.��}��$P��D��\����nQ�/�ͮ�������z7������{�gI
�'�8�7�[Rq��y~�����ue��M�����h?r�&����=%>xMN�l�G�����O��y	,��j�
�C^��lQ����:�+�Q^��Kv�	�&O�����u�������^�ϰ<AL�O�!shXIpԠ��֩=�ٚn���Zx�?��U|@�^`ݜ�[\c����[;X���m�	6��)�D+�D.	���7��XK_��"7���7����I�e��N�V��n��w%_e�d�
��'�r������H�������;���:�,�8�����3�=/��ڎ�f�T�2�1��h�'�[m�"j��a|��/�9�%�cu��s"��C3Q�t�)9.Um���7�b7���=E v����?%*�f���x&�`~$�����m�~Op�Į}b���G���Y�tP��Y?gQT��ӆ�~WjP �FN��c��X>X��zg�YT�0Ѧ��8�<�����"��e�c�*dK���!l)D���2%2�-�I� 7&��K�c6ZyOa�X(Ӹ��Z��[!��<�]x[S�^��Ae�<:�q�C��Ϛ�.�ޝ����:�ΒIZ5���m�c~���^�"U%h"?&��9ޝ3�:��*O{���7!r���?b%vB��X���XG��̠x�W�Ɨ<���L0���X
m��������q#؜��ڎ!#F��<��E��'�~�i"��,�����c8��}&�?���:��@\�	ۄJ6�����ƾ���XL�rw��Ov�o.����:Ɇ�3c�ט�Y� '��&�ӊd���vG@�����%���A����}��z��D%�<:.��c�`^�x� 1�)��7r���N5G6Z��(��ު	��V_q1�^�W7hgVY�&&���1�|kT�6�\�M��y* �G�a~��6�[Z�"G�rU��ؿDx(��b���Ԇ����:�+�i�m�x���ץ*��ܩ ��A�R��x��x����]0�_���H��~�1�.�?�/Rg�)�d@<7L�v<��\�ة�v5��w�s�)�?�̭��r�-�"ԪMָ���~�8��LPA�q�~�+���
d����[�'�do���o<�YR�����4)ۻX�N�;D�L�U�@D�Kb��f4��R�gG�\\��HPòkܥu6h^���o��"&ŷ7h��if��?v�`e#:3�Ꞟdہ�4�I����Q%YX�]���u��[�	�4-r�6�R-��q�Ѵ�D�j��-�����n�+��hi�>��]�r oMa��aJ^=���H��>f���-�>M+�[n�� ����� ����������"�;19���O��L'��t!]	�sd��43_��Z��[�G�,��u�#�8��m��0�&���SXI(��,5��Λ��X�Hqo�e�s���K}#j0C?#&��;4FMZ�0��[>g���*����n�,�{��b�KW3L-��z#�q�Z��U�݁����¼��Z��?_7҅Id�Q�-nV�������V��к7C�_:��:��Ҫf�A@��"�Q�$q 6��D��o��w��cv��݈�'��������Z�fX��+��M�n[.�C ��6�G��˾�b��pKZH�X��4�ĉ}~�l�%�o�ʰ��}ih�B�E��A�;O��9�^��T>��~ F*&����V�a�KxӦ�r����KV�E	[�
O��.7���/�s>FAs�d�Ǣ+D�R*?8�g�+�+���$Wx�V��-o����ۤ���,�d"�[of!\�HU�&MIe�s:LA�U'�w�4���U�IE��>��
S�н|P��ϝ,��1���髒�J��l5dX{�3�A#Y�>�/Av�Î��y^K,�n`{���&riy<��: >q�l�n�sH�
��qC� C�%g����'H��V��Ӏ9�W�*� �h3^�U��C�P� ����]1̃I��k��4�|3�8�!�m/�g�#.�Ot^Rr ��ꀯƗ�j+��$�1��F�6Ua�à�m��9"z>M�qe�����k�Ɣ&�c���;�k�Bf׾-qH��KBF�����R#7��
��&+��m��]��/��0�MJ����#�lkVS#�y3MY�^�Ik��"q}��Q���5��o�TwI@�p���O�������?7�>���clkOC,+���Z�-�J�n+Zn�Ms�����Ao#Q��HJz+�+w,&P��q�F"4X��kA�\S>��vT�sBWy"MH� {\,�ޏQh��3��P"�0M$�Z�"$����6 +Ilx�=�
ޕ��,�7�u��`I�P=�j��Q��0���h℩E�F�вZ�)�;��ͻ��V��c�B����Mf+��?�)b����B�O���/mbJ��^��(d3Iw�I��$�Ӻ���e�v�$������T�+�{�!�����R�2�`�=�|��� )��&0��
S���:a�l� /�2f#�+��z i�?VZ��y���5k��b��B˴1���΂+xq�k9Ό�w2�$�������a�� �t ��+g�t_o��C��I��"rmG��ĺ^���b��_�+��r���Hn'���x, C��"R1�n�xۿ��B&��w������>m��t bFm�����W�&����=JS��%�� ,�u�݌,���QR)��v���_io���.�A�B:t�oGʾ1W��r�J3�M��Ϭ�r=�h&5�Pv�`sbđ�:GHV��2QT�`{���4bf𳕺�}P7��7jk���
ܪ����k��D�D���"�w�����z��X7S@��������U&����1�PU�͙ЙJD��n�m"�~B���"���O4����z��+�����ް�yU~�,�f^B��xHfс^��*IM��Ig͚�+�Y�D���mbs<�E=��T����B�������yL�g��(�'[�+=�MU��DlZ݄��3y��B�R�a�f�4����YS��:'F�J���j��}3rbG|�f�5����@�8'�U֏�H���}��&I����/����p�!��8YMo���_��}���.K�V�wq1�y��9�3F�U	G�(����a��ϊm4�Z[#l�n��,|������y }r�lls�������%C̯y��K��堼�r�U�/;䞚%v��]_7]e���G6V��ҽ�f&�c��-�2����)X3��ֻ��#��yx�Dj+g��Ah�^�0
-b-�iJh:M]V����A뵶���M}�������[���na S��bRsDB8%k;�T��<�B^��%"YJ�S��[K&���~{���[�hV��L�ޞ�:�ǡ�Q�4.u/��WVC;�"r}�p���X��T$%6��ɗp��\ݵP~)�hڭJ��pg'(�E��{��Z~�6&�͔E�th8K��VZ!ܯf���/�E��k`G�Z��4K�?k*�w���_�90�}Im��OZ�5L���tq:ppq�;��0���d���Q��,�cׇ��"ҋ~�7����!#�hK�'�� 	U���L�GX���VwЁ�˟�S�g�n�)~h>�S� �E�YI��o|÷���݃_�z�\�K��M��u$c�G���:��s��L��HPf/!�l��7U\X��8d�o�o���I������A�dv�A(l��Z�S[i+�BFӎm��?�aE\�V�iųyz��k��8�1��y�h���eZ�U�V��c��i���д[���ǹt���t��j�;���r����B�H��vO�n�G}ٲ`�9�u4�jֆbs��R��8eNӔ���W[_I+25}|U�&����H���]/E(�'9Yq����� �ǧ=���Y�<ס�o��H���=�ww�.��M�ò����_i�5ӅG{��˿callgL�~��$�*�07�����6�n�LVM4@�Zwg�O���F���-��zݩe�Y�������)v����`a����ѹR�R��f	����k���'8{����*Ue�*�"@���ϛY ��]��W4�R|Xy$ֈs�����67ǋ�eiՠEm"bT�-w,E>c'j23���Ybr|4�`d�4�Lq�4�Pp#Hc��cjB?0y�!ueŁ��R�;s��b�:d�r��yb�&�~ ����ɡrC�۸�D���:O�k���֎�0O�����eE�aZ���U{ڬN����`7�D���&����q} UY�ڹ;b���e���"��%����N�ђk��싽��U��
_�^�"X�(���NZ�n)�qN�/���3%�D�T�@�����mo�b��d���!�TEh3x����0���Z�!���)�D���kx?�m�g�
&9�l�����G؝s�D-JL��
�M�y<e<ջ���L�@P1&*�IO�\�d�|f+�7ɜ�-��b�}B�e�KM�>B�l?R c�&0���l�Y��6����?ҍl�N���}Y� cH$�h��
j��}�j<S�Ӌ��<��5�HPbx����)�Us�� 3o��!˾o�g�ie�FM���^C���M2��r�i��I94�M>ӝdA��(ž�bY�8��)V��������޲������:<^��:6�g�@m�"v[�y�:��j�>��cZ�' �r�p$�y+QTA�x<9���x�M�_��?�
�%*����E��Lo�%�o�G0�S�G��wF�o�Wk�JəR��'$w�nS����XQ�Ȑ��0"i�wR��F�/mfnHA�!j=q��\�77���T��6���#�P����d��u�jϣ�JO@[s
�s�� #����Iº��=|eX2�(:�0�]�r�2T�0�00�F�<F���(Y�=U�K����=����o�AG+5'�Bo�fh����T�> (u��޳b`��m)X(��b �h>��w�d\�7k�T�6w�)��d�hӀN�
s�y\�����������W��X��h�B�y!�[�<�V��h^&��y�W�=�^�lJ��G�����n��vGln�9i�"zL#SR��Y=�t~����K2P�]�~0Q�吓u�"�����F�@��w�jO�[�l��!�ֈ�PACSf�zRy`Q0�3�E�7^Z�X�r�N����Ya��4]�ޤ7C�T�%��o��1��B-�]o��������&D(H_>��N_��׍4��-~Zӛ4:;�r3{�5L����'�:�q���
���P�r\ �$V[�y�c�Ċ5�}�9��=�[m3�=���&V�:�����B)�!��^��${���A?@L%�	 ���Uu2#8.ċ�zX��Je���ע�%Ú�$�vq��B�fkk���nҞ0V�\��Ka%�l�������6�ހ����qՀM��"�]���v���:t�*��!���^��>F�u[��nQ�'K;�;����U�!�����mo��}������q���%�ib�J!TqA�z�(�����D7¸0گ���;��Lp��˻��x���M]Xy;N�(Ͻ���Q&!�r������Ը3@�Sg��?_$�I�=�T۪˧F��##t���"U GY�Y��ʳ;9���90�&a��N�F�)�.�1�W����3��	�f�d�c#iAT�6�)���9���ǷD�el9JC;��F�w&����r?w���QB�F��"ݣ�Wƒ��~740�%����N�$+���_�q_<��Y��tF��"ro���|q�I8M��S�*.č溌�n�'�%�>y�A1�����)�$��c �^�1K�+[�(�K7ژM�?	H��cu������E�k�jC�	ϫ{�[!������H借��K�����n�i�x_l�>�����Ԙ�=n �׊L�Zo�*�Ì�>�L��rV��փc����A�����|�gڊE9�ݗ|�����οS��.�ev �>c��(�Ȓ����ז�r��Τ�y�Ê�\~� �,��6P,�G�?^�X���|�]|�!�-?�n-3�fh�M�Z�a�׳��q��w�/��D���5EMu#I�"lh&���5-Q���I=�7�Xp�F��Ƣ��E 랅��pl�K�թ������)ޯ��	�)npE�lڒ�5eA8��g7��� ��q8���Ff.���D�i�T1;V�_�T+?4S<�k=���d���C���ĪS{0#"�G� aK�y�����.(��}w��(S)�A��V4e�zedJ���r�4G���T�S9;i�n��!)��˞6V�DA�����r�����m~���?������xR�'�hS�Z�H�ў���J�vY���Ⱥ�9@���F<ǡ>��-�Ҭ^˂
<���qQ9���CE؛�@�H����h^����?�V��W��D��K�f��g71y�u4��} ����?}�e���N�=�vR /͝<U��IKKrs�
ȴ%�q���DշQ�=C�?V����wS8��<=S�Z"EEM}�3�
9H�0u)��0������z#S�d������^����Uh��[�wï2�&v�ux�Ӂ���:m-*0����ѱ7�HN�%s'����.'��Y�omu�ٻś13��0�5 7�t��Oۉa�MPj����(���T�w��:�Ia��	��`gQ��ړ���L���+~�	o)+��>K�vlw�Ɣ���H#gQ�E�}�Z1k<s+c�-}��S�����]�lG�_��Q�{ei���wN�r7l�U~���2�	-��:?��%A^1�
�����LU��:7:�i��쓌���p�^���a�$rPt����šF���u�8|��d7v�Į�!�"Զ�9^|�-�ȝ.����C�m������`}�&my�v���4��; �p죕*���TdD���:���]7��V��\fhsB��)��������vU��b��;<&>#��6�^�
�{�ԑg�lTC�ȁ��*/��� g<�7y`�J�Z �_1+�)0�T����Q�hO5���󫡗��!c�U��2&���ҷ�R����f�
�� �����
��nM�{m�J�*�����څ�O����R��(�-� C��� �Y�%�gٻ�^Xc�6&�U�7�GM�RGt9R�S�U�aũm���^y�����q�Z}�e>o���.��eMOBQy���{}��Ǹd�z�
�}�>�k�S��� ޝT��+Q��� �3��Vu+$���Qe�ϓ���fG�Ff(�%G�9�zs��@�^� ��+{���#b�$����:��r�9��
�0��Ӭ4FW��C$����=�dqZ�����|���:ըܻuP�n��_h\qk�"V��GG�#��.xQd=��ò%;���ozI�3�V�vd�]�����{�<A(C�c5Q)��$����b]��,:�~5]�q�;���H�#Ϧ1���l$�O��P6�S�
=�q���b#�<R�U�3�l�1��W�pcL�����͒qz[ڬ "��/"��N������$�Qѻ'q��m���֡!Y����'9� ؞�A3��%�S��-Hɽ�̈́S�1�_mAu��%�XYb��
�V�ݼ�v�P���Mt�-��-u<~w�L$�.W���X$�6Bvu���x����,�4EPCFV��?7�U�W'�.n�d/�d#�݊�6D��=����{o��ьS==��E��+��Ҵ��#n{�������d p<�N�gf��f�nzSD��pw4ÄzRGi�-B4�rC�	U<�W�u��/�K!w7�;_Z�PN}�)ф��H��,=�K����4�O�!ZS8�E��IZ�*�u|�ϳͧ�a֧�{N���KgjS�5	z�ݠ'w��k �Un��$EJ-]É-G��b�����7m|��F�p��-A�R�{
:��4@)]LK?<���!�� �6�-�!����ы�;�������u��'��5=9�K��U��5��2 ��5�'�kY�m��-�����7�B ˸���(��*,�k7�ª2d�@a�$�=�B�c�^(������h��������-�ɬ�Հa�����K(<E��lo�P�jw�di`��>�1b7��� ��W>����<�.ڦ}��4X�rk����t��#��0�<�\E�k�.p���nȊ�
�=�+ZO�ck�܉��*������D�$Y^�P���>�f��u����\̍�#��#]��.�_.k���{�"@���u�Z��L�+���TY��_�6���/ �����wS:q��&��Gũ�}�[/8CD)�RhU5���Bzȹ-�x����y�4����_����,�?;5Ȁl�"�,Q_sQ��'��ب-4�p
z�
�>P��K"���a�	K�>�u�R�F�h�Lg̀0~my���O�n%r�+S�i �������Ï[�w����I$����1��\Ƭ��Bb;/�g��/�RC�S ����n������%��*��> ���W���U�S: �'�g/!��x"�D�����۵��`(J1zX�&��Zj���cRK�1�Xz�8�i�q�=b+�A�륰�tC�%*K�	���\
���bȘ�$���@nuǱbn�5N�I�/7,.�����V��c|l��W�9yӦ�����Į n�{��G��"L�v�X�����Ҭ�Dq7}b��~\U�Y1Ϯ��X�������h"�[�vb��2�֟��7I�֛<o!��v��p���+5]Nc��</��k�1��:QvK�E���?�KT�F�0�B2&�[Ĭ�{f��\����\�pHݽ��R<M�eɲ�s{��Jh#z�b�my鿛]?'
�xNwRI�~���Z*�� �U�W4�.ݺ�Fv�h��:ۮ������b}�	M�&�U��]X��H�l��#~p���W�HI���Tn�fG�&���ܞ��M%��Q����p;�R�u��{�raD���V�Ṕ�,U4n�2�ri`�n��M���]�&�-` (�k6�^zV����T�3>�Z�N��lN�w�� !�v�&�!��&m�vrȀ�{������]!=��u�e�n������N����H�4��Ĭ��,�WNT��%@��Ds�� Z�^х��H}}ށ��M�~9~�٦����(��<�G������ۏ���������G�J���?'�|{���3ٝ�mCbz�>�G�f�[ k#�J�:����#�DK���V��'�{����Q����]@��#b�l�Tk��'�ul�ju;>O�T�u���Wr>YZ�^T�*$���ږ�ګ�/J��^p����4�4:2@�y�j,�#�hÅZ��ҧh�ļ?#�u�r���W��;M���W��3 ���8��uf�H�����,Y�o>y������+��uS_v��W<^" L���,�
���j,���S��<�+�T��7��Ag�+r�HNb�`i�]�*���>JL�J��=��I=���#�U3�1_�oW�Z7�$�� �jAhDL�W�b���6�VCjNwţJy?�t�G����H���
�p�!�W�qM��w�S��QC~�M��u�_�m���.pFj�&�f�=X<��@��������~R��jM�R[,���Q�+ȗ �7��a��cx9e	��;5L�'�=�[s��&��� �W����zX+�XE�R%)~WGNyá�F|g�R�;[��� �(56d0�i.�mp�W�/������RnG=���k��0����O�5��?��1s/�!���s���־��d�X+,/�x�H-"��XM�I� �]T;��=���ɘ9q�����`GX8ok�l�����Z>8V.�l�坓�b�)Ո������O���X`^T�N�eR���7O��9��n~�+՚$K�s�h��E0B���,�ꞵ\��8[0��5��=���R�
m�H��jge%"lo|hg1� ���f���4O����N��#ꆁ=d� PV�U�Z&*r�Hm[I�rѭ}qh��i�Bu�=#��
*ZN������1��ʢ����{��3`���idߋ�cOy��F3Rr>�:��s?w�w�`iI9�5�J}7��9�[Bm�'���$O&������Ԁ����,�9�G�1�wp���A\�AB�bL��ĸ�����@���'ȸ��9��v��<D�6� ~�>����TR��ER�6�+���bd��z��[���Y'�+�'HRa:iʴ�9��xx�:��gV�=lk�Vև�=�3�;�8.s}Ϊ�W!�L�NNT��k��ĐV$z#�za�K!�I�؄@�A�a_ݹ�MQ˫� u{��/M���=uN4���O*黐*����������=��I�&��L����a�]��uT�dC�_�-�l�F�
g�����'�+�ډ5B̫n��I����r���F�����cFz`ψB��OXʗ���/AL�5��9����T��-�Ʒ�l��ί��-�<��M��|D�G;
�
�5��+�$����c���i�������vB�):����F������|��ڲ}=��c���*����1o�[��o1�3��\E؜أ,o�R�H�A{��{��nR�c��ã�@'�+����m�<:\�TV2��ֈ��b�L"<J���zl��?��9N��kL����D���Џ�Wz�hn�2i4���Ca�5�$�Y�ܱ��xw�L�s._K\-�
G���:E	����׸��X�G;��A�N��rΟ7<��� �8�b�I��Ox!��3~]5Eҕ���1���J7��yJ<�iU�J$d��Iv)A8�'oLԜg槀�n�)3�n$�y+4Эq:����&�5�;��<��[��ゐ��Yh{(�S�X�7�F<��fH����I��+\���9����1����/Ũ3�.[vtW�q����[VB?�o�"��͈������?(��E�	�Xe�~��G>J��9���GE��h���&
��9��&�
���F��L�U�L�tΕx6P[���ljK	�������ԋ��z[��i���km��ҏ��|�^+TPa�%y�>R�]����~<��5�=�R��*>��g8��0Z�I�j�Z:[P�_D��S���"2� e:IOr%�I9�F��(��7��`NG"��-� =�;;�i[�}F��3�8�C�01َ��b�t��5��&�C�ۅF\�����sb&��x8�:^�!x[	��e�[Y&*k[���Ƙ�6�S�^C�R]�`LIo�z�	9 ���0�B���j��72�p�p#Ҿ�����&����r���������%4����)���-��B���Kx�v�;/�<ߒ�T'K���<����O��_â��o~kd������#�M��E�j~�l���O3=s��<�X�慚�[�1҆'����hF����SR�Ki�}� 1+�k��,�B�y��dY��d�N����]\T��p����a���}qN͜-�2�UT�ֶeU�JǣB!�I�+���Ag�'�����Q���b�E��q�r��	��"�0�Ԁ�����<�o#�Q����_���<~��a2�n0���*ρ�9T���i��u������=rj�Pp�x$h�S.W�\�v�z�T[�%���!ѽ/��&��L4�Ds< _�;wsb �8�/j)6���Osǂs�!8ޙ�p��h{�܀���篁	H��1���3 <[r�e�/��'�~���K�����U�CI�iF�8 ���)r%D�)"�o���H@3�<��$�>��CH�Ԙ@r��;�������~F_o�]� C�v��<�P�fiŮ�/�\��3�p�Y��c���a	��>e�x�b�2���-&}n���s��'Qcv]�~k_W���U	QG�7j-H@�o��J �{2�����H?L0M6�'�3�~~̗ı\�Z�-�$f��n�|S���&q�k.� �?���N�^r�(I^��'�̳k�_ݪ�o�����n�U�gqY�1+�&�i\��,���R�P�-{z��Ş�a}�C1~�Mui`�Y�:Ҷ��u��Vy�u@�����)jR ����gV�j���[��i'� ��-'Z5�c��/K�n�j?��Ӭu�E۝6\G_\�?�L�䧘�_d�Y`n2������~OgP��T��w>�[��D�[b<P=0��
���F�̴яեX�Ĳ��Tr�~N1�s
�@^��Y�4��R��𹆵����4Bz�۔��\5��{6?Z2��4�X�x���.M@]S���E��m#Me5?��oz�f��,�{�,�N�qs�Va4f�	��oL�% �~4mCF9�h�g	�r��څ�]���v*���nG�5")�����(�?�N���5JC�h��UĀ$�(��9m%�|(%�9�R����N�����c��nlVal��M�XXN.�L ;�QvO��K�v<XP����Ni)@W�غE�-%�%D����x��"�A� �����=c�q�9���z�@���˓a����-ȯ��r�p^XV"3�#W������%m��}���,vɺ����b�Vr#�o���:g�Λ�l)ˣ��H�R��ҳ�'��I�M�߀�DӸ�S6��nX&#��E�t'o�|TW\l`?8�m�ۜ�� q(2lW��gl�W�C|eY��&�Ѷ�.�A��r��`���.SHH��}007D.W������yF��KT/#�I��������Te�,x��~N�޲>����׊:_�!���Kce3j�ڎ=H媿���Q�0�D��P�,?;����`�ٹ���B�u-%@��7�x��}�&�0v	 b�ni�_�9��у?h�1�p���u��zʤ������Z\ 1�@ª3NB<�T�J0��<]���(�=�b��b	m����־�I�f�,��W��$�^"�u�z����G�~�ީ��wc�t�ǌ�tsS'G>�*�<����6�߈�_�I�C��Z�î2��6j��Ŧ�h��㍼�@���ڄ�dR �ϫ��Ο��t�,�ZD�P�i��7�Ϻm�=n��l޽� ļ�n�fR�Uz{P!�͆��OLc LCQ�ί=�>�����A��������%��A>Z�E����T��E89�U�z�h��O�Ukі�o���Oꔹ�->j��N����jC�ȉ--�=Á`��w]�z���mQN�7����1�A�5Q���k�:���nՖ{	 �%87��4ET�$|f��A�G��{a�gɹ=�xĀt@��O�[?�tߔAKG�BP�s�F+ҧ[c$��6O�B`��ۄ1������h@���$���h*��8��J�șѝ����>��+�P��B�@�$�!= K]q���l�t	��ѿ����v�v�ӳ�xe�:�]��R��D��	�V�]�Ҿ�&֊}��4H��:ڰX]V��5Z�������
�,��w�;�+>��-k+z�/S���κw"m�I��f@}���,�Z㤦 m�2�-w�F�H�ߥ���-*�n�=ҽ��r�;c�|b��+g�9x���k�T�Č�����[^[���� g9fg-��=?��^v>��6̕�-�6�0��؉
���YI_-���� G��s�iv%)o�s>�r�t$S;����Y�_Z���$y��Q�x'Φ�\p�0�G�Q��w�N�V	�J���|�4���tK��c�\R��s�$"�'�t9���f�ȭ��Y#eQ5�lv񷊻�׋�,��<��Ǖs$�{�����UX~n珅�e�[�L�rR����ؼ{�=����if`��(�#�>"��I$������>��'s�k�ѱOx1�V��]��$���\�o�6����uz�"�����dWI���D-�嫝Y���9=�J����W��Yt�8<=.�B �,�����/}�P�_��$�@��.1ЁvwՊ2^��Xj�I��i�_B��G�vV+#�1��d� �������8q�� \cA��r�_�6�χ�و�=�,?`�V��F�Vꠍe�+�L�T�X����܄k|�e���ԑ.9�Ip����b���3-�4���.�_��^�D� FJ2��G<�t�?G��-������hQ�>��O݀�4�%�.���f�PDF
+J��и��Q�V�{���|=b%Y�C �0�Zt���%A���F㣛�fR�����$��C�q~��V#�F��ެ����ʌ+_�3[�&0n�d3ڶeր���i`����+eM	���r�� �����N[���^]�he6�p�JYFK�;�Fv@\��Y�P8�,T1+e眼����S"=��(w(I&lp=S*j�L��H�@�,SB�	�y��l��
0��*^�A�u�}RdtU��0�{rۇq�Q���=���t�C�l������+�\���Z�"�Jo@�+Y�+�V��]�:8��Z֌y�j�V�3�	�R�@ܿr�h8�<��<��#0����ò��#u��[Be�k~�p�,-��>��B��a�f�/[��RY+9�F�dw��$M�4�.��M�!´��Y�%*�e���3ޝg���V�s�M`�0��8e�g)���,���B��ơ��0h��L����o�@`���?o�R/D�h컵O�6��*~8%w���xB���3�2C�ܡ��ȡ��o�mG~�e;����#@��|���gb	��$��S�&���ƌiw�r�ly���OC�Cvq^�Y˲�4s��n�U��>�Ε��.XNf��4 �7j�xf&+�}�ja�-�d�6��c8�N�UC�vq	�auO/O'����[�m��-}?a�!��-N;�ɿ&�k��s���t���ޑ(����t�i^ѓjhX��:b�U�l�gz�SH� ��Z���R��S��z�#�a&5�$�t��+��n�1�Zmef�Ԥ\��*����+n+��
�r]!�Q����6n1���5�	�U�A݇� �ϼh�h�#I�On�tVi��3�~l���P��m�s<���씇�gs�1�U%%�i��u�{ڪ$oy�<�9�����r3��Qm�D��}ӯh�-z�.�,��~6���(�OT��Up9U�;� X2�/tM���oߠ3�R����H^(�Iӌb��tG;���F�}�T�Г��43N�Gq+����������ȭ�$g(O���z�Rl�m.���ZZz�&k�J�5Ђ�5�Kk��߅E>dqD��W��_��sQ��d�|�2p�ؐ�����xEz}A�`�	F�"T����x���1�����>�>S:ӧ&w:�`�bGT�~����C�%���{�?ˬU��7�F�UQ��,���0wx4?�m�C�����g@/�%��ة�zNk�R�!wPj���iB�'/D���n)�ϙ�c�_��.�>"��*��M奥��7O���}̂w���C��p׈�>�Y	Sv�i�ACψ��������5j��(Cp��Q������~g�$�Xn��~j2��I�e�g��F�e�{yD�0�$�1�F_�JM/}:�JӠ���Q7���ۜ�uA7���k�9z;�6-V�7fGp�ڜIcS�-@v��pNWǸ����a�B%�r9 �"C|���QH8��L�=5�:��`����F��oDv�򓦥��3_�EB�����������e��������'R��S�Fpb�<�y3�j
޹~�4�c���Ϩ�<ElO�l���U�,T�#v���4t���H��##V��'�z��c��=����7�'2w�n�},܂��S	�h�f�CB�|��!��[B��X ��D���!��m��=�a�L��3��#�#�@�?�B�X�n�k�G��k�_GN��K�'a����#<�H�ՊQ��M5�������N��R8)����ƥ�k��nM�m��٘#l�]�f��ăӖnQ4˛lJe.�M%����߻ޕ��z/3 �Yg�`��]ˤ�i�����$���1_���cC�
��?�l�" �:�Q�P��0���UU�ڇ�5��N�hA��*�c�?o�WF��C�>P�9�k��#(F��H'��n!S���h�� �w�P��=���:�ٔ��,���MTM�S�-�Z��
��td�1�T�Vw�[7l�b�Qc{�.�Y烖08ǱDu�K�mԤF���ߞ(l��I�fi6��@�潾�Hi�?6��a�.���誴@=�����倳Y��"wMR�tuJ0c�����PD&
����)#�m�H�0#��C�M!��7�@��&P�/���}a񠧸u�$�u���'^�]�>�!!��hk*�|Q:9�����<jy�b�q�.���S�-� ���d~dd��:�*%d�G:FhŠ�̓���ߪw߲[cf' d�|�V�T��Ag�C���d�|�/�ԉ�I���X�O�3�'��0fm[�����C�˘�Q�^�`�;���L�3��������+����۲:�N�l�|�|��MF�#�N����.#T*<�J�.�nU2z?'<~�m�X��6���M�di����6�v���Y�����d�i�K�B͚"L7�����ylWi�[\���.-,q��%��l�fn���n���0S�D0#�k�Ŗ���{�ɻ	���(��&���7�K��m�/dm����Gd�g����f�n����%��b��>��a����4M�G��-����j�>�ְ� ս�#>.j�&�I��߿:����[�6���c����z���ʩ1���"9	x�$���@L����BO�!4P<o-"&����UL3���z�a�f+AD|lM܉�}N��o�b(��e�&N��%�������)�kl�h���b��^���@�����(SV"}���qH�4=��'S@ЏY8�gz����׳�\��O�l�"�o������#���RE+��䪥��|��v���?���#GU�t&뀴���ܚ��"�b�~���R��E��_1Kf���1[`ͦ�dL^i2-dU����ꔍa.�1����'{Dp��U,��	�!4�pV	�|��S=���C9��h�~<�zP�C��,`�m��=�s�����K���i`��B���p9�V-�9ݯtYJ���~�� Ꙧ ��k���|/��qC�P���Q��8U#��peB2�Кޣ�����;��(�����P-��0U#T+m��ݢ��mo�(���\w�u����k*���^�5)�`��dщ!�f,G��y�V&$�氩zS5䀝����8�Q&����f��U�+��Z��{����?g'+ZCNX��N�֬����q�g7�m'�t���X� S�a�~�Y���A��*��������.!�9�<bl��'������=)8��_�E�ǣ#;a���]f����A�u�y���¦���'u��LT�����[���|��b�"򽀰���\��	����$/��p���4��˽,"�����(EC��7s��ˤ�A�w&Z�r��r%j�PD<�tV������
�qF'-^�r�A*��I�瀞wU�(�ۊ֍@�ҋ�=!(���&�[� c�\���ڲ�LG���$KG��G[f<�]�O�_��1�M��|ez�e�fi��˜!� fS-3R�\1��8�v����x�d�2��.�p@�M� �殕�?
���Ԇ	����5��W�\w�P�����.�u7�m:yv�P��fA_Ү�v��m�#{�~�S	@#NcIe�W��d%3.b(�~�G����)��T<��
��*��hh����Ө���9kWN���^���F[!i��WE��
j_D�|����W�s��f n���H�Dfc��С�`	��� ��JQ�B�����m� NJ���m�Xw��sUI�=w��-9��� �[�� Bc����'��id|`7ۅ�I��_���1L�뒦ѿWX���N��ݏ��l�h�H�e��u<� �c�MZ&�+6F�ap��y�4H"�:��N�xڴ�IWÀ�h�v�'h�.��(%l9�t�Ga�k)�NtB���w�c�ڞ�L���PʯG���+��s(�^8p�m�$�z�dS��S�E쓷̗D ��U���J���Gc�1����9r�PB��Ƈ!YOa�s��=�����MYU��X�.�x�c��EycN������l�Z
��n���������R)�3D�~��7��[@�?�
����\��R�LF�Z�X���cgK�6?I��ّ
�wTA*'�(��s��=�3��	�TU̩t=5�u�b�Q�z�n`/m�
�P$���)�#�;�����`�o��'�S\��
2��I�R�Vd~~�"�c���[q"��~$#�&|߷�dЙԑ�i���������:��Ш��sY�ݱ�̔�u��!i�s�Ӵ�_@Y��GUm�u#���v���V�|�&@ %��!vM�/mi\{{�+�j�c�Ϭv�9����k>�2?~qHT&�	���ݎ�=�Ŕ�]�}���	=���3]&�/_�t�8��\������(���h�*�P��A�����%4���$�4I�RuX�毓t�[hs���'�x��u�s������$շ����.#n�����]�R��}��X�x<������4���$��c��H(�0����㮩Fv���]� F_�p�=��L6P�<|%q�ۼ֠�ezZ�8������mV�ĥӔM��<��7z����J!L���X��ɾ}���j�@��ϰ�/�}S��n\8aǂ� ["4�hk�Y.1b�0hyD}���M�u�u{O9N��ivx�����L�h7�IT�<����s 	c%��#�4��(�ߴF��9bs�������>��I/Jvb-�*u�׉T
�!�e"����#D��&�Qu#�n�����Ĳ�V�D����ª�If�ye.��[�%J�<z2�~LYʱ_7�h�z�$y�3������Ҍ�RY�(�n+q�顇�f��5�</IT�B]n��f�{�;h��[Vk2�R�?͚KS�ņy�2;xƅ�r�-����^Q�'� S\8/��mlWt�x�?�rΡ�/�+�ڃ�$�~o]��h���lB녆=�k�+hX�n��k��;��L��7w���f��������F��eCf�\<E��ʩWJ&�p��1g=D ɴ-@-�)2b����&$�PtR	���.��4[���I;_���W2:N0�~���SA�(�w�O�GD�����)MR�z��c���+�^���Vm	I:s�2�Γ汅��x�=�Qi��8��fHen�ֶ4SA�ܲ�j�`&�$I*^���f��vAE��6���{�/�z�ҴEg=��;�V�7��ЗN�=�o��D��J���7���&��������\6�uA2��k
<3�heM��q����$���i�*IM���_����,� $�:R�A����o�+��la,� �j4\�m-p���kզ�"}NQ3U��L3��C�O�#�,��7k����rj�Pd��PZ!����T1�t����>�j��l����zo�r'qkR���s\�ܽ����/�̩Qx�;�߬�_���Ȑ��-� w��j����;^�.s�n��3-��L��s���p���G�J|�Qm*�XӋ�O_;�"e�N�If��մ_g(O��>M�R�Ζ~m�1�7��#(�	f���SYL��,��@dV�����n�KU�R#Q�,������&��.�\��@�����0���L�������>(zXh����^=�<����(����������$�?�b�SqRԢ#�F��uO�-���M�>�����Q�;�����?Jh6-F�{(�&�MOpM�:�u4��U �Y���+���C7}�R{4{����UgI[m���F���+E/��7Q��Y�$�x�;��GxX�TQB�V0�m�d����%*�5�wu�J>q�QrE5�e���$�X�n;@�YX'�Xη������!mn@�'B�uֶ�c\�� 7�O1h�����?{�%��V�A(���E~�h�q1P
Z��M%AA��	.dU�y�r��H���i�%:�6W~u;oi�حB(�^��2៭��e���>�2��4~���qD�8���)n�m�#k�J�ש�|��A_�x�x|��_{sB в�k�y��P���I�����,踝���g�U�?Uso��T��_�J����+Q�ʅ6Ͽh�KAW�)^m�� #6q
��^1���Ia���PR*M/�W�]ly<�\)��"V�f��q,��&g����+#�OL\���ds�)���{<u�� u�ƃ�N��GMI�\�$_���r���㧁�9ґ|LW�昈۲�N�zx��%�s��ĩ@̱{ŷ�&��S+�ʢ	���d�$D��h��hLs��i�M���[��Tɕ�n���A�8������(:�oS���%z�z�r�����3����#�:�n���'<M;����?�(��'��$�8 �0�h遝P�R3�� ��N>��q�t3�N�\% �UJ�deeF2����&V�B�6�mF�^�(�C�
��
�I͔IT@�4}e_���0�Ye1�os|�#yg�z���ٛ��@��9v�M�jZ�bnT�L��Bb�����v"9F��� ��J[�3�,#p2���VN�6�e̋<K���.$`
C�+z���W��DkA�" �����-z׉9��C��e���DZoQ��ԩ��+OIG]W�ơ��,���A�Q&(H���2�^����[w)���Gcx��c�n�X6/=��|`0��xXmӢ�ӟ��,���-����s�R�O�l@�g|5	&��<�ck��B����'����$}̼ؽѬ�&M{�, �NwShHmh�>Y������M��B��ZY�����͘�U��s�%z�n��4N����9G��(�<	��3��τ�M�w(�e�vy�q�x+r�:X��V����C_���?`q
��F��smza�'Wy��}����U��K��@	��'e�@�VA��#m��G��e��s e��Ut��!U��Ԇ�M�V��ɔ���hw�9qn��3�U�z&���Nj�z1���T��<W6	(��#DX�U����������4c��<sW�IW���C���I	��{=���"<����ɰ�N��͔J���m��d����b�P�z����r1�+�h�-��6�� x@��+���C��2h"����*}�YMD�R�c��k��4�+���wxde�*�B;�ꖑvأ������V����W
�xy�20�'�����{��&g7�6�⼸�֩�"ä�>bȨ�B|��gF��-ʲp%z���\n|E+��U�'�����N�hq}�~��^���@�D>�/�C(���Eưf��1�	M��6+#�}'���8�w ���(�ٻ��R�WXۊ��ԍ�Ĉ�9������Pt��`�C^/O������_w"_D�y�,"���TK�Y���7A��cЂ�lK��R�	�~;1`�ݻV�|��YA��HH����%tla2Θ��4���dD�s�����k�}�m�g���5�5#D�C*ȷi�����u�� :;�F�}[��g4���mudi�H-�c�4�iz1���̦',;G�pO��f<�����81����q"�7���p�`�P�j݌rPr��!���*x�g�Ǧ$���������~�A�����NU���
 .�y�t;��^��#蛢��T!:����h[���VA ����Q��aќ�c�G��d4������"vnl��k�o��U�W�w���y�|���U����E+��POO�'����!�7B�[�]��y�Ey7�sD$�BA�<t�Y0�ęl\`�A0QQ	�N�
�ɐ��T.HH��޵��J��|k҅|f[��}��X�qW�*0�R_'���/ ��i��g�oc2�i��zz7�K��a�A��.����(9��N]�P�L���i�ʹ�Æ^@"H�eڻ�nF���r(�J������j�E��� ,I��7s�����f��Q]�T�Q�}��k(�����"[�G�-�徉9�_Ç��;�򑞥vH��/0��}V�醥�/w7b%q�ϻC��Ǘ�/s:U��~��~X�-�&'Ԏ�b�G�nFw��O���y���6�/;b���p���l��m�q�h�݀�܅����l�+��:h
���>}[�'����[>`���(�y:�7MM�̦/}1_�DXKZ�vrO>�Re�2�v�#��w+�ot[�N~])�;��������c�V��p8�!���cJ#S;z��M�l�	e3�ڮ��(&�=Դ�GmȖ2;��q�V��S	���ِ�͂���Z��4��J�+K�;�Kp�}2���M�+U�k��FI��$"�"L�xb�xr`/N���8�VI%r�ATeW�}�k���$zEnȽ�GD����X��!pȰ�-W_,�!�Z��l$�(J�� +}�ħe���x�ts�����S��6hd&�R���E7���o�2�.�z���km�);xK�]�_�����zϲ�Z�MJrSj� ���*A�4� %4��µ-�44'[�T	�
�������T��-�`�|'�m�]�T���#�Ǫ��Zp(m�C�!�����tA��9>dظ+/��PF��ToJ\���-C\�w�+'Z������x��x�!#45:Ls�����b0A�U�M��W�D�Od��y�,���}��7��9.G�m��?aXNb�xM&�i�߆7��>���e5�)��!��&l�O����$�DG�"sg��d"Lk�E�=�HR9]H����!�Cݶ����i���P!&�!�-0A�=�yU)��u�{c�Ĩi��R�����V�!&�Y��tt������J�V�[Eʸ���j���٭���Ȭu����aG�IY�����T&��s`�,Z���C�G��'�g͆���#V�z1�Y�� HĸF�����rQ���u\N�}S���5=F�!��4�x��i�ܰW�>����@`yvĝq��S�K���&9��˹e�0w}Q.��M)fj���3�v1�����I���4,u	j]�
�;S�n:S��D\d��E�6��,=�������7�օ�������|/��©C[��U뵭���l�-�@�l�C�1C��ʁ����+~�dО�Dh{����n�B�+��-R@.��a����Ǿ{�͹� 5۫���\���<8'����0�K2rӘ�����!j�Nc�� fpV�H�E�hn]���1���d������6���b��zCߔ)q3�-���[H��Bv^��b�So@��[��_���(a��qϕ��1�%����혱���� 9T3��&�j>���Hg�e���j}	&58<8q R��\q��ضi��Y#,sHN!�L61xw=���G��)vs�Q��KR��{���M�&��u=��!r$�Ԛ�J�fM�=���r�g������S��JK��S̙Z� �*�+��T�b�d�$��p��cqe����x��ė⧮?e�=T[�])� �@z �!�i`��4���a�q�p7���5�X^U �F6�s2��e�v��Xj�X��}�|��R;�ϪQ�d�gj�F{W/u;�:ta�^8F�U��U�J7���3淍#v���n�ʃ�	����k1��rǐ|�E�ᘇ��,S;��֪g��<8�D������-�ҩԈ_��spa�L�F���>�2�n�������oM�km����!� ��~^;r�tא�F9��L�ޠc-G> ��A�|O��Rv�s�&�[$�u q8^2����ic�*2;d^o�p�(�&{���l��C�z�ɧP8��2����nXM����_&�Ȳ|���莯��n�� 9=z���7Vx����|p9�+�WQ����9[N�vϓ8	�	��ao!��z�l��<��Mk������M9%�_Y��?'��'k~7;zD,M�߹5��~NW-�ECm;�u2���{/�]�9��3��R���{����[�lK��l�~Z)�p�>��1>c(����|V@�m�9��(��"�9Қ�r�M�/��C�$��I��Xd�Z"���ET�F;��7�ܤﭧ�w�Á��nh��9���y7�%"�Y���|�zD0�y�U������2hc�ۤ��(�L�np������O^J����� ���Ly��oZ���{��h9&j6Z�
�h�a�J�^��@��N%�Ѷޮ'�R"�h�h��Imv��j���dL.���rb��aM��Ѹ�cg"�/;%C�a��@0t�}VAu�v��N�&��{�=[4U��ĥ��$eQO�N�V�݄P<k��/g��&S^���ۀ�A���	����&a�V\fnl�����Z�����b(KB2?�Q���
�6D��Y4�H�4�Q�}����hx7��D������^(4)�4��P@s	WP�qu>��:�7��rBd8G�����w��7*��[���3�G"�e�ʘOޒ޼���\���(Q����1W�  ~��]�
��.�7�]���Kؾ:�K&rV(tT-?@tv3�0�L�+V�a��"T׻}���$~^3Tn�4� �^��uN����"��V�T�9��De�U�ɉu�P:��nh��d\R����j]7��k9oo�fJC��˕�u��*��Tgy�t#�13Q�`���6GS��w�'�<�}�5޺q�V�b���D/�����\g��޽l����b�s�쇀�Jcd9��䳒<����o.0-ﯖ}Ŵ���%Շ�W��� ��+R���P�0�� ! J��λ�����2�)}~��ϚC[�~~֨)�? ����e��(����(ĕ�M�z�z���+�i��*��*�Ɂ!�iC��(:�kZ�Sx�x�sb��A���/n]��r�u0Eyf�]������.�,��/o֠.���EԦw�:a�V��N��8�PF�>Lq�LT�D�78�qČ�\�AAA��蜖���2��CjN�N�`K�x��r�-�ņ��ٱ�;��0>���	��j�3�r�K�~)[G��P~Uܴ�-�ڑ�Kゖ��$4� �k׾K~�.�~O�v S��ꦩ-3�'�!��k��`+I�ч=���ԃ]�GCV��"����n:Ȋ��Lnj������=�\
?c�|i['H-��I��hk�<�:kw�kb6��3� ��ym��~e�f0�kV|RB�����|3/�e�Mv��,g�f�4�D0Ҭ*
\\oI�1@Z��iz�z��5¶�&���B2#ˉs��� b�m�������~�T�p�{���y�L�N.�MIij� ��B���w����E�SV5UUn/X�Qt%i�Gj������w��������/ҥ�<�qH���6����h�
O���P���h�E[(�0�Y�ʠl1��eV�?v������4�6�4�#b��ϱ�8��@��|�{�<�	�V�;n�W����,W�I�����i1	,�c~�Ț޲@��(@ȉ��X�נ�����ʹ?C�-p� ���!�a���p�%��;k}B��\\p"G�R�O��+�.���	>
h�����-�CVTC�fJI(�
6��jVF4�Sm6�~��Y��[\�F 3�CG��\�kǀݓ\�9eP���j��[�+����������������O�+���/���1�z������yԢIu����X��D<M���bG � c��ݲ��E��>Mi���!V��m:p���:^��b\f�yc�P�T׋:�qP���I����s����l����x*DX�eke���;,�w��cY�i�Yf4�[<��,n��ʘ�k�	^�g��^���� �l����J擈����D�Ѵ��0��I��"h�X�2{8tc�@*/���.�.�{��t��U��.�w����G�A���(��5̙~K�=z�{E�@4��jP��Y9�Sv���P�y�*���}��?����Ü��p&ұ(yO���W���=�K�xld�U}�S�v�\��B#��M��y�����tV�����D��60>���6w5(~}���5|�,����E%����=�l�d����"͉ox�/���$ 
v�R�#2V�P��o�_�f�)֫�
@Ǘ�A��}�k��1t�.ڹ�r�ґ}�!�H6v�6P�_-���E�Q����!���g�B��-gR��1��/
�o	�m����0E-���Ƙ�(G�z�D"�$����¶��߹�j|�@��hz��q{*l�-5��
!M<
�l|.�YZ���Yh���q����܀ �TiA�,׷�|�^�H�2�2�JŃ� i\= 4��9�f2u�Щ��zl]���~M��n�=�"��}P}6��9��M]Lm-�*^��ΐ�Ɯ���bYa���[�S��/��a�v�9��Τ�쵄��O�I�]�H��N�N�?ᑟ$=j�o�����Ɲ&�Nxr�����Z�M#�>R
��F+f����h�K��]+@6��qt ZIW�d�in5�.�M	���=���˛�W��!'���ù��]HX�'�jQ�WH���M�dі���K���&��Srz���Q�I�9%��;A&Av2x?�Q��O/��}j]�íA�q!=w���]�oFjV��~��)��Y���fA�h�Ȥi}�B�:?�� ���~g��+ߝ�;wJ��VK��U�f"�f&#,S���8@mJv��T����C)�4�������%�Q�w1SU@d�z�@]
��������3�Z8�8#JҮ��c�3��u|���ἑ�`��>�ơ6e'Lɏ*�N��Z����[8�b�'&%y�wO����|�GJ���θ����ٰ�e�/�c�Lc8ym��f^΍��� 8��d��tJFh���\}��{s)�������ec�>��H�%�U�`<�p�n7�Z��V��{O~q�2ڟ�1K+�4Ww � '�H�;������Ӷ	2M@p�7�q��2fֳe���p~6���u���R��B�x�C�J���2�pG�l��V�D�͗�$'�s���@�?U,lo`�	n��\�K���ݧ�"�|l���͍-�^}��<�p��Y���,�i"����B7be�]mi:�W+f�"�ӝz{q�<B��칮����Fr1Ƭyol��L��R2�+뗧	[�5ꠓK�aT�{5���0-7_����*Bm9�'��_����5Ʉ�|����5�w2�ږ�������m�IJ���.N{ �]f�9.`x�e3;����Z$�B�n�$�r�f�_��j;/��*��q�yǇm��b���6�)��݇r4�;"/;;�!�0��H���H�5��Ef	�Qg�O�+z��OO�/|n$�����7�/ �����St��+?&�5����^��'��Q��W�1?kA�V���>֏�G7�B9�Iݣ�����Z:Yo�4�Y��O��K3*BY��M�R���߫�\=f�M�2 oif�],* �\��/îp�p�����FÄ���<@�����������'�D�4�ys��!�}�����S$��߈�*�z�B'P��l�ؘ�{k+���c�9e�᛹�o�V�C^��D�=�O&��鋾�� 3�1�\�(/�s(T�D�b�\��-L��@Ԝ�s�x�)X����~-k�r�r�0�p���i��|�0��-�"�G�y6Ӿ�x{HP��'!�O���[p����O�T��&/�'�T����΁I�Qu�B|� (�J�y��#���5�a��*�U�/�0���� �K�˦�~*0��%͐������D�R�ܧ�� ���K �o����3y�0%~�g�G5ۅ�����&�_yhG�>P,Ĝ'���h/Lu�m����R�}a����PS�U�����y��@5eMG�A����C�ܯ���p��M��ߥ���̧֕�$�D��m�oi#���v�[���,E�F7I��:�:���V���l#a��m�V���ˎ���r�h�ϨZX��h����Y1]�\,T��V�{�& �<��:V��x�X���b�`����z����o�����*�]Z���oo抦�S$�H�y�j[8_l����Q�}}��u�O�R\<d�@"������P:0R���⦟i��umTkUrCK	�$h��<�C��G����l�r�7��43��"j�7��j��,՗&ú�-5�8�bHȼ��@�[|L�~?\��(X�G��1I��C�ό�˗��P�������a��L�j��(�9c+�KN��9}u��1m�T3W[Xv��,�5|qsw�BI���h��ۥh��<y�����Lv��J�� ���հ��f��NR���=C{<��@4�S)	_uPnِ�d����E��$ǧ���w �nݖY��Ͽs�4h�e��j�] �A��\��ܬ tL���6�Դ娔i8ƚ�'��#@'b<��>�B�H9��s�8Q�h��:)��!�����U�Bh����q��������������D����C��}W�D%��R��d/�/n�Ee�4[[���f[�5�S��v~@ǂ���^���%�3+brV�G��_g^��x 쮯_��;���$��2����!��YBЏ���&���~�kP�j�ƃ&F!��Q��
ta��I땚���M�K\�e�)[��P3W���퀻+v��mk]z������9�X��r��k9)e��nRP"b&r�$�YO����"�-��(�9��ܗR&�k�d���e���b�	!��פ�wN��r�G��U)��x����ܒ�ljd�R7(:M��U�#ex4eF�"�=j.��b�*�b	~mϲ�WX���[~�f�\�7�ܼ��m5�,(WQ�a��34��.J|�9z�Iq�0"�6��í��Չ"����p7n|�	�<���)o��'�lk~"�35������BH��/�K�[9W-�W��3ݯ���fZN�ى��b`@��ܨ�����F�(p��d^1�ϟ5:hG��0	���_^>��t��ez��YJ'v���M�����KĬ�#��'��ED���^�g_�d'0�a���t�+�h��]�π��#�s�D����T�=k�uvH���Rp�f�'�x���ʘ�s�f���������D�r25ܙOw�?KKFv��S'C��Ws2�G{u𡘿�����R��B�5�.�9����&�h�K)����_2����p��R �6ޟ��_=����&�x+�L�jw��tn,�b�I��J`��[LA�j��t?��Jڧ��2ӷ���pw�2�|�{
�0���I~�R�����{���+c����ܞ�4L���7�2����p���'B<�rC��C�����(����yP�`�l�u�C�.�c|]\0 �r*vo�P)L:�v~���Xh��Q�׆Ў�U�j�Wh��?m����l��\1ѐaˁ����Ey����{�V苮8冺G3�SPa��V�]s�&�����ȅ@Q �z�u&��n���Q�ǢuaZ8Q��?�a�u�Rf����!K`�S��}�*.��H&z�2�W�7k��*S/��}��f	�4�ӛY�U�΅��\�~"�	�j�R1H�}�ӡrkYP'�9�>�.�,׿�'.�Ғ���N�~���(H��yw��D� �f�����ֿe�O��׊��Yu� ��Y|�F��̵Qw��H�_�6�!��>�k�\!�#8b`�.�eP�?�Y^��4_Ob���-��{�ӏ��f������f� C�.�s��^�܅GH���	{e3}�}������hB���0nD�[�����Р�kE�r{x�<(�K 6E��(��}�`Y�y5�	\�2^��゛]F��3D�4��KA����[��_8�� ��[�0��%�L�jJ����t_ŗ���������%yŖ���bB3���v�o)?�T��]so�uI�K����[��\��M����c�	��G��0�T%��K�zH̲�V��F����R���{�nn����{��^Y�,?�����#�iwrqo�V@����O�BZ��[I}~��yK��Y9�ީ�׸n�Q�l���|�OM�Y''���5������Z� 3��e�9'�>��(R�g7u���4��d�|K��Q\��ae:{��J�IdB�(�kŁY�6$TD_dȿΣ�����9�U�ԝMh���ڷ$�+j	����kh�4��~�)>��4u���+�r-;�U����2
$[�&��}ד����w��"R1 ��вu����N&w���>�O��p����E+#g�˥8 g������	~b~�"��JO,"�_�&E���r�3&�D%؇� f6��1�y�h֪߿�Q�k�_n�;,�6�c�x04��ߣ�7�E>�B���T}���Z�o���@��F:3s����)E�juj�c�u@�ȧ��We��r�c�v���V�����Rn��zV��Ы�\˨җ͢�9��pf�l�':�Tk��ߜ�0��KC�:�l4��f��9����i�R���\�覗�J�h�N街$!}��P��w�� K�0���HQ�+������`�~��Ծ�汍,ZȲ��kZۺ�%�l��������idǽ��(�>�JTͼN�ۄ�����JDQ��$��Ќ�.�qU !���UGr�H�&��1ޭ` �, ,TA�#3�1�n�{:��,������\
�h�3#9芈���|��r�$^�YuXtyY1oҔ�q���,�c���v}5�^X<�9xX[�E>?cy�c�?F��R*�K����������0}��N/�fa�F��SV�B+sg� 0f�g���2̌8i${�W,�Y}�u�FD!?h�0u�O&�/�$Y*#^@��X��o�����[P����B��� ^&௶�jr&Ƌ ���h�� �\``�ܦ�r(���.��M���_޶e�U��r��1����^�m��B�qE�$q	���3�=���f��O"]�^�ZP�r�p��g����7��H�P:`8�� ɽ9�e�$�^K�R��@#��߱"0��K(�P�����
���iE�1b{�<�[�)�L8=v�@�+O�B_�y]V�c(��R���x��w1�~VB��i+���V�!�P�lɆ� @�3����s�~	r�P���[�&$�ԊA������� ����q����(lDw���1Q
F%#�JL�w����0c�%�lҙшp����6ZUy�����C�7�*�����a �
!���)���Σg��]�`���)�-_G{��~�uD�~�^�E�jվ�]��!�s-aکH�"�g�Vi$D]��"��U�e^^As��Ev�Q,o	�/��,��yr��L��ܻ6�w�,1�UP+�}
&��n��d6rk��7��Fe�M[d�M���	n��I9�}��Ұ���>�(wD�H��'~��΀���B���9]��S��}�w���VM���q��r���+LI�\�� ���=m��j94ĺ�9�tɢX-6�u��D櫯C)���Y"7Xf�*��1��xn>���^�M�q!s��g>hȷ�#/�!@���w�SOt��aB�(fI��?Wg���_�~/m&m �4

�$c������!՝���!�{}��z-��d�3$�,��q9V�#��O�G�[ԩ.��c�TI�鑟���v�1W]B�jLbp	����o�$�Z���=�����uO1���×�cȲa�c�O-
��Ȕ��j�f�h���)P���9�u�a���d����srh^dG�i��6��e�y���$P�����~���o,'�-��v�wh��C�#����(�8��/`=�8��)u�SC�W�N�����~A�L8��3�vӀ=���
���F�E�TI&~��%�gg7�kl�[�?U/_�"Q��>dM�hs���uPUH6lt�>��U�j��J�M}��Uf���١��B��U�i��&�AA��g���㜁šʄT�[�7T���u��"���2V���Hmc!�2lf��1�e�o�J���{����n��"��y����w|������l��>ߒ46I��	QԆ��˞"B� �*�J5F���~��G��@\�ݚJ��ZY~q��Z�M�EBC&>x`p��O�+FX&)���B�
]��t3\hW��A5��1�!��~�%�'o��%x��j�4zpl��Kya=��k��b5��Ys+����KB=���J�8$�j��|�%�Bx_��ط8M�IB��%����D�t�Q�\�]�?���c,4�v�� ��(T{�5�vQ��űǨ$�p�t��>r�ဃ��A�'�7�'/j�ţX�hf��U���n����(��ŀ1�+��'�
N�mG^	��^g�+۱������)a|��
@����
�/,������9A���K}�� Kg����S�!�C�k�0rDP)�m[2��K:[�ӖU[�˾Bzi��5��L9Eo��z
ׅ.E
��{�����:�Ӗ1�mp[��X�( 0�,�`����9�@n�s]ϧOK}���3�~/t��I���6m�`'��!��ZR�p�hͣ���߽�  �钂���oy�<O�;�?m�y�4ޮkP:�(	�L%� �Z�=��M+Ị�O�_j�X���h!��'hˋ�a�~�07{�_"�#��2��z�f-T�cC�hU@�Z&�YE��j�eW��τj܍����D�I����*���"�ud���9���g���~j��.]�]���ѴX�2��˵���ǽL�x<i���Q���$Ar��@b$B�U��K�L�����7�[��2L�`L9Ͷ΂��]W�G��B�o�G�!�#�20.�kP�RŦ������4MA΃�J0�l9��a�!P�,�:�v��T�@��|��,�V���'
����	`%R��u5ɴ�6�\��|A<ܟ��΂ݐ&f��wm&0F≵Ġ�a�1�e��q����L���W�ǌ�㞦�2��~���ӯ���b��C��w*��ɖ�;]��\���O�.!B�ԇ���� '*�D�/|%�M� w.o�ݘ�A���l!l�&-��M���~��J�<X����FZ�2!-cH/�{)��u��4���?e���m#U�訥gAE�@����ޞ*b�Q)�#
�����O<�5��l�.���ϧ����=���}9PA���� XQiF��R46��d�A86�MlZ#�m�.��OY��ғi��zf�Q7���ٻw$��/#������>��']G�͊��s`�My�ϮG]:��r1�U(SʙO&��*�򛀮K&#��;O��(�W�q�G�߾��7sY������cZSu�o5��?{/�I��!J��?���!��j�Zaۇ\Z����y0Y�w
h}����h��Z4v�G�֞��~��Ut�׎�-�g-�(*���Ф6�t���P�,̹Z�_@���c<�\8�6��òම�[qt��4��pa-�h"Grv-�.4��Qu�� {4U`�냸�2:�H��w�K��!o'jB��א�����GtO+b�jܯ�.v�?>��mQK��X��p�F�� �L^�4��Ƶ������m`A����͟w�����!���Z|�F���;�bFDt��lkf��Y�R���~eQ�u�������.���A-aI9|l�N����pc
�~8�o��M5�4d!�#�1�N�I!�._=�^t�"�(_��@��1�J�|V�
����k�x9;v]ߘ�����^7�"c�>'�fonZ;=����'I����.!�F���n���������b�Rt�htgO�Wi�f;)���8�C=0���N:�N�Oo"���R���7����
p&y�UP�<Y�]j�j�D�oi�`D]���l~����
	�hAt�0�����V$���PB�Cꮏ$FQ���~w��8��uQ��f �>�q5��0�P�_�"(s.N/��)#��/��7�ϫ���3�>P�2�F=�#���Y��S�?�a�t����|b��2/}Ӵ�A�C�q������R����w�P�S.V�y�G�fn��ss��`�=�9G��(�d���hDA�^��Y��E� {��٩Cƌ��5·~(D��Oc��:�C�<�'Q���͔�w���ͤ�$��p�(�%&�?���?�&q�:�<�h�x��0� R�C��\2�;�m-|�S��Q�EX=��Yc:�y�l�
4@�=$�	�yW�l�%��L;�I(wMo/k�m��J��G �f7B'AK�B`	�[����9��K/�P����*��+�S�<��g��^�|@������wj����x�o~��������3)E�w7]�BN�܅������_)�a�������/A�#i5m�j�s/�<ӓ5>N}D#�&%��w����\�'�I�&����5;v3Hbm'��
�Z����:�ñ�ɸ]�S�V���\`$@�%�uQ(-lB��_�BNG�d�.�H
�6�@�id�U]�p�wNߞ��d�T)|�0X�ԛ���N���}�L��d����R�m����n	��C,2!��`��)�����U\$2׾@�V�������~Aڭ��:���o �X.`�h�h�f��;���3M��)]&:���U�8����Pd�?�~T��(�������b��Mֻ�)�g.!?�h�'�s�m��k��KK�)�X�P�g��Ґ�JBC�P��� �u�Dx=�ݴ[�'ЄhP�l����������1��r���FZQ6����]o��������,q��W8�5�o��h}ҟ�|�4�F]q�G*-4���L2���,�g!���=�aĥ).�B؍��fW-2�4^�೮�iT�`w��W.���lp�E��1F(���DE{CR�1xU^a�pOsge/�<��������{l+�s�U�>O4����c�rmA�TJ�'J9�x��u���7�zY���(uuQ❲nt	������m��;�C+	�5Jy"�$樘�Ĭ�W
�?���z����BY���
t�%����Hj'��N�
����G��r"#��P!�虷
q ��y�
@��b���p��]:���]�j1�z&KP�UzKL�Ef����	�Ey�	짹��Lz�-Mz�����F��%c~�\K�]5%^Vݲ�j�H��j��T�4�U�6S�em�	�{6v��H��J{� 9��I3��YT���`eFv�.��ұB��x����s���ɷw�b�}U�i)�n��������u)k�(�\$�tȔ_�r|sPjT���������L�ur�b�;'5\�{�Bx�~*���L5:O�A�i`N�3ueZ�k��h ��'W��?H��������M����"V���t�d���-v�g�@{�� f�)�A�lV�XȊ�� 39�YS���w�Q�I�ƛ�h�t���0{6�U�i�����`��	�<9�'P����tC��%ȶ�H��V�#�7��� ����ę3��D����{_�SNr0�I��v��NIP4�e%��"�RUD�C�zI+�{�N0E� ���QǜGv�E���a�5: �c�Ҧ1:�ޚ9mZ�`Z����#uM,Jk��S���f
9@�6�!�w�r�5�tOg�𴍷=�UH�/u�g���N���jك��(.	p2T�bq}��w �����.�wsq9�ui��r���N��?���^@SFv���P$N�u��C�ѹ�B��K�����tҨ)=���P)��{��l��^'w���a���!h% �8�'�sc�10٨���`~w�8,�� (��OѲ���\�q%R-JQ9\H]!}��$r�A��VA7�U]U�$�z-{�$�C���cѡ��a:�'��<i6�_u��ɰ#����I�p(�	$C1ݜ��#�Fv��et'�L�����Q�Z/
�!]� 8���;b,u���7�筽?���nn;�%?��"�=皣w�e^�Q=k��`��թN�9ĝ�D�p�NR̵�D�K�O*U���Ib-�X�2p�8q�M��0a>�?x�.�%iZ,�r3C����@��CW�#���>�s!����}�:<�����{����� ��}�H�����+w�j��Kv��2�Mv(�ޅ��|xz��_}�yg�;j����ҙy�yD L��+�O����*� ��T��/��jS��>��G�6~0Dxw�&�0*A)J�	��85D#pt17�Z�J墑�݁�Im�w ��* ��5��)}8�"� 5��]��������6;
��ٳ����}��L�DSE��u�ǁ��|ƶ-E�Gi�c��T7��.�~���t�e©�0~��k�%$A;ϣ��j�X|D�rԤdn�p�4	M��@����!V�V��0 (���mln��/�&�`�`S��+�U� \l� 7;s-�z4�׵���o�d��2\������9����X�֤j;�a�o���9XT$�uYMDȍ�N]�g}^b�_��V��̍�\hgL�V��L���I~��� ��E����$&<9�I��9� �<�r�������3�_���g�9��ޡ!�4z�w6��ͥ�J�4}��b٧r��Ô��"_�2��r�=@�|�e���2�=**v ��!��G���*�!�����Y!��~o0�Y*&^�[�Ku�S�J/ݕ.;!���<TbJ����M\[�V�qQ ��}q�������u�� D���V1��p���&P����)���\�ܳ-H���|�!S�~X��=��h��~'p�̃�'��vˀL�0����®�#��K�U�4��J�H{�gDG��sR��q\��|N<Ԃ]0��/+��J?UJ��%�j}`e-/����J�Q�����|b�4�sGh�QH�h8 �X�L~� _������Q�q����F�?�No9��V�,P���N�N�QU�GxʪG(S �c����(�ե���S��U[�ΰ������Dꑢ�7�B��JӢ��rr�R�Lw������%$h�MmâN��%��R�+��9^��A���������NԆ�K?g�B��gt�� �{�����[��V���l<��,Q4zW)
<ԉ��4�$�=r����>�]����}ha0�5!�� m��#��'�+
fϋ�_}���Ց����޶����:��ۉ��U7���th��3ŷ�\����!u0�Ѡ�pd�;�d����sC��0=���H�k^��	ިv��<f��:��P-�4'c��$t��	$�4��W�PϢ�"�i�����H��v?8r��sF���	��y�Yx�N- �U�ݱc-���=Ր�L�V;P_��`��Ttގ��#�7��Ǥ�i[,��y���,��x&�����#2d������K�HA줼�M���M����ǞLVN�n�k�������7<�l>��3<q�9�	W��;[��}�{����&�F����-�.��g,��r-`��@�v������]d��p��BE�O�Mj�iO�9 ��ү���u�2:�Um�Z��s[n�N��L0`��n�ֱ�n�����dH�;O��1�`�r��
�&1�my�������8��P�$�J�#�[pY"��xy�����<J���(}����f_z�KW�fG���b3�V�1��ePF��	�x��ҥ�(�䐸fA��z�7�K�F�SfoE]�����W,�ӥ��("�1�T��W��/�O��K���{�L��X�V0B���R�c�+J�j��:#�$��p�g5���5���gx�����AX�a�Kb�8tʀl�V�'���I8�ޚ@BO+���唏����<)Zΐf��c�����:���]����\�ɗ�� Bv���yO���	Z˭K�C�O�5sr|;Π�([��/��'K*���$7f2��u�ڼd�NE!Dڟ����)��|� yQ���Ț�F<�����7�@�F��(Ͱc����̌�H�F��ґ�H�:��I����B�����(�F@/�0����K7��/�f�o'2��^�Zd�tZ�t�\�a�yH�Q���&?y����!�����yZ�g3��)Co�3��X��^Yϑ[zɵY ��K2z��+h�Q�/u֏<Y9��	���v�H�d��h)����r�6���څ�_��Y����G�%�vo�i�Y��~^��>g��5�6*Az�Ib�����]���0&ַ���O�l߈,������Ek����۶,���/� \���_�0p��Nb".��*q�&P��9�FuO�j%=�H�EZ�b����c���o��7��0݇�R��ymٸ�o�X0��F%{��{�Q�d��MdÐ�{C�D������|�%"��
4�Z��g�Ɍ�72�O�`�A�y�B+/hoߗ��B��ǋЯ��P�\�ܟM%;���{@i��7Zv��p�8�ʷ���؉��;�t�WK��D��Ru�I(���*�����-���;�e�^���K�����)����_�D�Q	�b�հ�T*�o��� ��n�OD)0�8j�ɶ�M�e.�-p%7�"�����F1�?�R�LL����q2J��V1���Z@���t�UN����V�g����{6��&�xs_�3��n����i����h�>�2;��z.i�^؄�޵�Qq���\I�Wۋ�;K�~(�A���i1���5�`�Z��φ��
H�./+S;� |���x�hJ�3�y��VY0_���{������֛PF��I���+Ű��(bH��pYfF@�z�i��dΥK-&G�ɣ ຄ�JV'% EɌ���$Jҹ�o���ހ��V���2�(��[�e���;B�l�) �y?a��/֌'W2�c~-d���[_�M@��կp��S�&�-�H1��%��,*�"oWq�@P��\�W��?��h��ɰ�0����`��ĸ:��7+�����E6M)���$��Dh��օ��$�/�"�	�7:�2Z���_�c��z�}q��1)�����R�)��^�����7:L�O��� k;(���2��ϓ�;P��V�tKRs����U��~��w.���U�"�G�|����?FUo2u}���u�nK�#u��Ш3,>��<�����%�Y6��\|�^(�DS �QcϚ3/�A(��C �ɃH����a��'(����w{�0�n~ Y$'�t���68{Ɗ�M~���MCi=wC�`�;�P8s�	DZ:�n,�r���zPgZE�%�EE|mق��@s�v)X���u-O����vc��H�eX��Ȝp,��b�@Ki����u����l� 2A��a�:$����z.mE��9 ��&R	,�ܬ�b��si���tmF�(�9���@۲�������f���z!��|�e����t��Y�m��9�HC	RVB<f��:s��2��u���Ò#�2ȡ�O7X��Ig%�t;&����\p��;���8�	���ٱP|0NݪR7m�DZq� (����������J4>�̡��$V����U�@E5!Y%���ƺ���[�މ���i�TE�Ф�AtU��f؝�2�/T.F��"xv��Rk���$�Ī�L��=�������d�]����
�@h������ۅF ��lj��r�@y쯇ۿ_���n���wF���盛:�MMc�;��+%@v��j��(#���N:�b���Ū�$�0�r�?p������q;x��&@h�cYƆM�k�3�m��r��DE���<��?י��B�ן��Wi��?օ�L�����!�|��na(=2��>b���wj��Z�i��j�A��M9�T�A���υ"�W����V���:��޼#�_�N����ay��Jjh�z�7ʙ�#0ǂL�#irz����*�لs����P���=E!|��jJ�>D�Ӆ�ϑ�� �2� �)����Q�7�����Ihs����{��pf���#��#
I�^�Ο&�2�"�{����:��mze�N��x|V�ݫ'�G5ټ_>��oau�vs��_��NǨޅ����2hw��oe�<f�J���	�z�a��0�d�5ٗF�\��---Mˍ�qW��E��a�����p��X�H�oE�M$c���R�2�Y��7\\7t /��Q�Q��D��A�ӊ�c+`Trgq�����%g ��pv8`��I4�=ҡe�(9�)6�p
*r>���]�_�����Lқ{�����T'TIB��ԅ�F��ƌS^-��`B�?<�1{�Y��)5)��H>�~��wB��)^G~1�'��P�p��z슔	��2��p/wB��|[��D±�k�U)�%�R;'f�ue��*�~��=��4��ܠ\�����cś���	�� ���cuק��X_ӛ�l����Т:z�4
�Ao>$*#��{�V,ٍ�#Ɉ�R�g {a�ҫ�zW~?��1�OsH]�BT=aUb� ��T�?�h�Y{p��5Wj
���C ���o� �Z��na���ӭO�"���� O�T�f�q�C?	я9�ʰ�Þ]��z��g�Z�`1bp�&�|Lz���$}��<��l[�QpV�WB��&�c��iϙ�p~ͣ6��ብ��'�O�����Ǳ�bSඕ�Z\"J��� �2��#c%����5.Ɓ�.\�g̶������S�Qt���)=��ܹO[��qم4�,��k�n��o٣�q�@ߙ~"���� �Q���_!Zf\	���o}�-��9p뙦�G1�6��- 0X�I;�?bo#@�
�C�8��]�d�1�)�Op���;��J������: f�`���Q��:k��lǕ��iH>���@9Q:�{J܌I�����D�o��u!�+�=7�Nj�7P&��lE¤%��č�dm�pgꫥp���l	���-e�e<{.�nE��T,���ӏ�C�s�������y�,�J��2R��/��b�G��2�6�Y5�0a��&,;͵Ƞ�&�69FH&���>��o4ܭ���k�*���*Im)�M��f�)�bףJ��~^v�-��ru���3���`4����ךئ?� CY�lh����UVH���������h��	��f0���Ա�p�Q~#dx����]TGx�� �5���i�#�!�j]���Av�ӮY�v{��A�<�G��T?���"��9+]�"��GT�k�xO�ǭ8���u���������􅴋�����kYV��`�<eP�ʙ�F7C<�H����l�ȴ�;��)��!x�w�\ﳠ��$�S�=�7���%+�;:��7�X*�m6G�1O�E�$�.�LԄ�gW0�,� ���8 s��k�d���4�W;M�:X�ңM����WFM�eǮp���w�[-����;�պ\�Z��l�u�/0.�-i����dn��!��~G������O�L���LN��29�k�Ţau�*L�Ar�k��8<m��g5S-ʪ}e�#�@�cD�JE���"\U�M���5>Z{a*~�h6������<^U�W�?
b�ck��{��`Ij��o�TJ��z+bB9��곩��=�]oU��u~���I6��ߥ4J*Pt��K���F�Wܣ�?�V�����@E��&�PI�6^ �]1�\��M�oSH�b�W���<����c��Qf�0��#���o����,���~e���&�*K0��5��u,����B���\�Z�6��|D�C5]�_ĥU��v���Ԣ�e'�Jw��7gq�'}h��7\}��O�Ղ�D8�*�;{dg���T��Y"�i�J����5e��XJ�.�j�-��%0�;�:�&=goz�E�D'_P:���5?��e�F)�#��\9����ʫ��Vr�M������q���W5ǲ�<��yr;}G�8(�/�����'�"L �Y����3_�b��*/�o�͢��َ+v5��R�#�{ON�=����d=���M^g1t.&{�Q;26y��MH<��p6�-���F�&���r�TM$$�6alv&$�>k�g|��+��H]�D�QM�h�ki��a�������4��c�nY����s%�+>#Ξ�+�7�ڀ�N0���sj@�p}.I8j�E�/?���=>��{�c�0����
��O��1�٭h�B���%Z�H\3���V�q�U4,�R/�k��-�RJ��	����h	�'5td���q�{����K=�ȒH���.���'�/�[j�)ط�Q%�&�yR"
��ś�P�%�3)ۦV��V0�w+�M�����L�6�� ��s/�����pX]Q�.A�*�N㍾�	��9��9�_E:�r]�[�A9�����-B�g�Ն7��_z�),0�`��#lC"2�]mH��n&�[A�r+F��H��ڍFc-=��9����`�8��x5A%d�X��lH���!�����[��(*�L�4Ĉ�0��#��b�;�^*�4̷!f����72��V�������u��C�b<��Am;�-C�0��w��̇Fz��ǝmq�䈯u�M���AiҎb�ꭏaM��dZ�sQ�ߓ9�!�b�����ySjp����T���X�!7m�>ťR��Wf��h<(�ҷ<�
���H���&UϢ��������
�3�ش��O��q����>��ۃŗ
S��?p��W0R�?��^ͪ���+��%~EkK!=|����m��.9��,���o���ڮ���$J_o����	$��|�I���Lƨ�$lcX�
*�<W��z� xޝS6zz��9�9�Kg!֒�ƹ�Z��uU#Dy��1.v9c�?7���&\��,Y�RtLa�j�w�{����%C_9L��bE��."����try䢥�$�>����Hʝ\�c�ϥ��|��X�j�d��/�Wn�|z��Q��(�a[��Z�t6 kN4�;��D6~˧,��t��`��z�"�ᤅ�VBkI��+e��{>��}
4�a����Vc�v[���^�})��U�y�
��I��iY���J`[M�-N��R���",�n �<`M�k9�A�5ے<��?I}�r6��Pdt��jC���E/Vt��2�MŒ�_�ǿ���2�2���o	܃�� 7����#FQ���	ʞY�$e�ͮ �m,�R!�4�C�9)�;f�O�n��R�vB]��DR��)�n��D�.�����<ܮ������_�����ҍ^���Y��7P��:�}���ү�Y.i�~GP#k勪[� �U��T�LFї�N�b�>��~�5���A��]Z=���{RT��;��"��������������TA���%ޤ��M�Lw�u��o�d�'�����7g.�%�z�Xa�`��4�_�;n��k�g��X��j��z��c"����H6O�H�7E�)����,K7�+췐�m���\���>%��п<�~5�u�/��kv��.���\<$�#�; _�ˮ|®�Y���vl��⎃:�$\������쥳Z�;�弜�9�Q֟`R���LK�c+9vU�X��>����ӳ�Lj+d?�x��>���^7��މ`b�h�������z���j M�S�I��L��L�W%~B6�O�����k�����Y�Q����b8��è`u�h�`��aNXNu@�>��o�"0�J�k<;<�@��TX��~ ��@ƺT`z`�m� i2�W+��+�>��a8�	��df5��m�f�&�̓��v��$�ު�C]��7�Z}�ׅ!�
��%�e i��juăŨ#u��0
%$�=���}�E�s�C�-���^��w���~ρδ��>�َ�w�wU���1�ٹ���s=�2>|����ëF-�'l~�9K/3�����SsM�~$y�>b�47)u�:5o'�R
���o8�P/
�r��ZeN��\D,my9$�Ã]wR�{k�G�x���v�#�j�>d��9��>5uzW37�W�rF��W[Z��ٍ�Bwc6����0� �K�X!���{�h�L�LU&�shvx����1t�h6�����à�Zm%�/<����gj��Nz`�{�;iA����:���w�yA�z�*N��W� �5�5�QL�]����w���6�m$��[���wF��J����S#����׉���5�g?��a	��
d��ֆ*K�z�㷦�ك�$6�w�l�-[iJK�rY�fb���;]9��,�zD�l{����m�bl֏N����(QڪSjȲ�p
#�vY�W+�gv)O�I�?s��1��A;[0��Jp!�7)G��1I
�p�����azS��oxtn!Zv7>5(��u�� �,����p�5�L����r�D�rv����P�<��=Y����`��J���-nVEz@*W��5bZ�F2���Ǉ'��ã��zz[�$(���]\Q���x�Þ9�y�h챹��Z�uĞ�a���a�������ʫ�4I �`�`L��>V.Tn'a��o*~o�h���7�S�Q<[
�u�(�u ��,�wV //�RYJq��ر:�BS��i9���7�v�?:�7)��-�S���x�p�61%n8�ӁF�-���Mcs^��(X��\�w�:�V�r���1X^��VXv~��Ż�A�j�P(�5�������Ke5��H�G���˻�ī����+�i�]�A�v���,�7���/����M���۳v)1����j\�
'W?���U�;R[̱�(V�⯬�_G�3�`���Tܝ��BnU0�Q]��I�%�x
��k;�Ts�Ey}��;7���)�&�{`���z5��۸�f �v G��C�o	�O!!x�Cӆ�6�"����Y",fpZrf���]8�L�4���$UH�0���I�`��#z�����d�X����ب��w[$1ޢB���������/�p�H���	��epP&�p���j�3R�M$�2ҥJ���:D��D5��}{Ϝ�s/����H�A��CO��[F������0�����K��~H��2�B�ٛX{�]7�i���&�Z��͵�7?��Ş�����8\(�\�#�������Y��m�,��Pv4L�u�Xo���i�Ҿ���Y�ٽ��٦˶���(JTҼ��wx-��
��"�����4��Iꆵ'�����D*�?W�֋��LM^+=08{D��h�{��0g�r9cb����� ����D�R�>��'�6�Bٜ���%��/��c�����c�����e�"�ҷ�6�����zP8AdĒL�I���AT�o,U��yżb��3���'>��BA��Gz�[����i�5��0�%Rv������|	�$�8U�ך�qr��fm��Ǒq4⫍�Qä}[*������}�1��ڒ�A��!�{A���\]d4�kP��.���ڢ/=�).��V5.ut])HCnd���4\P�I��#����K�����,^�EU�E)P�W3��E�ko��]�iK���Y`�]o�ww�_d�ĀgL���2H�Ѽj���R�GgYTI>�%��/���,�]�2F��?��mY��/��N��;{��=���r�����T<�o}�=�p^W9S���!)�IU���1�,x����G!ɖ���܇ׁ{ ��&�?�m���qmK��@��P�{�L�$%�^�^1��J�����f����LUY1��[7#�]g,ݥ/�]m��D$�St��]��.)<p�ߓsRM�-�ؙ��W��]�:�A��Q�mp#�����n*5O�h2� YD���}�~w��w����>F����U�{�D'�Yo�;W�ԮI_Y:8���@-v�V]DK��o���M����e7���ڒ*Q�W< E�I���[L�)lN2�%�|�F;� ��H�+b0�ٞ���F8��Zʂd�Yq���	��x��!f �a�qA���KU��[O��0�B��t��'ٔ�J���ld���W���M��V���bi����������e���O!���0ɨ�ު�VVQ�3��'�.�ZMe�)EN��}�#N[7G�C)ƶ!s�߂�m��PP���.����jbI��uYQqj\Ɍ��s�u�W�攱�
�sG%g��H��i3拾6�.D8Rɕ)�#HT���{Z��f�����
~v�}��[ �ho�u#U�� ��S� H�ɷ13`����lP���ւ{!���I�U�l�s�]i�y$�ǱF��!�o'ދ��xX��|x��h8X�\�:�Ep 1\�`����h���E:G_N>���wr��D��w�F~b��%�F�!�c�J$�zTW�en6{eJ�,y�+����B1r8a��י	��+�vZE���wf�u��tP�`��HC���J�����|:���V��;˵�ߴ�<��		�.V:s��n9;ή���O�L�g)e��&�����*u"ľ����Ɵ-���ka�ۂūbxK�[��FT�>)���M�uh"�1�VM	�q/ZSM8A��ю
�+��������C��Hǈ�4�|�cԆ6�.�%Pf��+=*��4�HZ1�W�ݾ�z8���i��Ou��7ft��X�
��B�&`�-�ݒ�1�X�K�C�����@h
oY�/�p�C��ϵmu��h,�4$�3[�U1��"o��]59`�	����'.��$�����`r����l��T�9�`���T��0Jp�D�w�����:7������L���7�{����i9	�=%eA;"�����W�"]�T�.H�P;�\ھ�B�t�H9�˅&����]g���b��滣���|K�&	]ҥ9~BX�Kq6����0�SQ��jG.��
8lG�)>w<��/Z�1R�y��o�K�A�7��t~KXރ!�@کG����A$�&q�����;Đ�`���!�)�<f�M�Ь-����%%��e+)AR�6�J�ԓݹh�lp�G ���{��+)��|Q+��} ^�ڙVr�/��H5����@H⣎��c�����#��R�a���}���@%���^����O&g�:�Uߦ��|��	�0kg�����rO�-�/dn}\,t"ISN�A�0��ĕ�)&�S^U�|�[(P���_K}�4�TG'JT� xVjN	�x1�����[���I��F���f�>��X�����|q��1(N\�^A�(A�a��	�(�hÌ� Y�i� �	����0��譛{���}�z�CBP8B#�ð��_�s�@��F44��E�J}�E��OY���o� ���xc��4�������fu,D��{p������k�ͫ��o!�йVT�e���	Bչ?o�ݘ��yzZ���H�ʌ��6F]h����R�����}.�&8P�}�(�l�NGzϞEf�%��o�E�bǿP/WQ�'��^m��o{X�B"j?coo�{i���vNkߨV-6�	��q$�[��|����1*�5���h�U���?�P�^����)�{���I��=[�p��9�Je�������F*u�Y�����g�S��2|�c�������<S;|/<
�΃G̃�o��C�t�^m\�q��\sV��4���٠E�ǒzA�7"QR��������P^Z�t��;K�ntޯ�Q�<p�3W��*��ds����}Y�F]U�7����7�0�#�[�k�{2(I�D�SE��m��.ʗɈ)%����ay��t�ҹo����������Fh��w�)�I�-}��qv{ܛb�0�-т%턍g�72ջ��zNjizt��k�Ų�@CE�P�e�c)�O�*�r����$�N�P�a�×y��ݿ|�>m
���c~6[Rs��H�KO[�%R��'��i.�vϤf��k�+��dF�#D��OmJ�/�	���Є>L��<\��0wB��l�p�.��u���z��q���&�-#\�ˁ�@��75~�17�� qZRΜ�b(Ğ-�ʰ
�D� ;𵪒AcRr��ܶ�e��G^��!��o�O�#,.䯗��e�x���'�������WȠ�4P�.�2,�������
�,~���N2ЧcBc%� �%��D.7|6�����0(U�U��ň���0�aцŊ)�� ���~��F :�����|����88X�'�Q��6cd�0Z<�45��z�C�]���S%N�{&GoP�� ��.�e��R6�f���W�$�4^
��K�#([!��n>zL�y⛷��Yg��5	�<��]�60?:m�]�:�v�ho���B-����%��Jr�x�66����>�ɫ�`�El���wl�1//sN��ٙpD!��r���kYy�f�[ő!P:t����]��߅@_O'W�z+{��G�
���[ |� j}��J���|����f���65�����X��1T�ʏ'͸�-8�n��"sw�&-ҏE�1�ʐ�:ٻE�w�Zs��5_HZ��#U,�y�<V�j�m�1�{e/��1uh_��!Fd��?� f)\��m��M8ė��).���6�HNzA\�y�׊@�reu�M${�{P(�l��^�TY� y=�5�gq����v��(��@i�L��w�$��)�W�M�;@�p�q�v��,ag
}+��YpeE짦p$��1�X4!<�	�ǵs+��ؖ[8�8�iwx�Gˌ1���6������Z��N\u���y]˲��Q7�9G� C�u6�>^QD��\�����i̮�,7:-�8��#j��xXF�]�ݔ�v��gB���X%�����#�P���3b���ʥ�v=ш��[7��]r�!{�s�YZ9���Z�? e{�-ӎ��_9џFH��;<�x+����Bj��%v�vю�P��3� ���aeѿ�b>�����{�x��O��1�PtKr��%N��нo�N�2���z�Ӄ��+�M ݔ��=�y3a�/<��X�	���>���,��j��ËqQ��92��D�9P ߰�3��e�	5�
����m\�m��;�Ͱ����ۺ�6�e�&h�K�Y ��\T(Ӑ� �V`�h=��ۖ�"�}��Q�٧L��S�AN��(8��k�C8��񋫗��{��.�w�+�F��m�����g�����@�d�q��%�����)�B��{8���N[��%( R����ڄ�n��)�)Y�\6�=�C-�+=���z(K?�겝=��l�<]�st�J��dG�͈��W�z7<B��UZӑ`�f��7������C)Sf�~�E�i|�3�і����K�F�,��]�?8�oJ�Gq階ǀ2�����q� M���sO1�gS4�����'�z�,�s?�@(�M���P�n�1|�'x�����rf2Y���"ؽ��S@#�V�)��Qѥ�5�C�55�vw��S��P��^���3��)�j[ M;�J�#/4jeb��5�·|��`\���qz�k9�le���F��OB��>��:h�Ka��#�k��҆���*���rC�7>mw����n��%]��
\z@��0W�z�M���@M6��j$�K�0��`���@�"K�~av�(�6jZ���5k��igO�j�V~��ޜ�~�.q���T*}��O�� A3�<[(�硆�ǧI�u�7W�Wa�` �h���ԉ��]���m�w0\#b��m[�oZ�@7�c����PS���#��d/5
�����TY��Ļ/����Gi-���G�������=�@j�� Xi������mZ�g���q�����xO�y��ߤ��R���m(u;�߾{]�ˆ��,I�~7�yOK��1q���z�u�`e�l��H���sמA��l,�_��������NCm�l�����S�E�ǻ�ՆbS44��,<���\p|��ى�����H�k�{�F{��}���T=ҸI�xqW���v(��W��>���q	s�כ;A^�ha	e�n��c�j�~�\�'�;�U��~� נ�N�[��@�z>I1�#W�R��3�j��-���b�Цq�飻H</<�T�*q�L2 ���ø4-�)}��~�����v�V�S��<ghP*<Q
R�*���e�nd��ŏ���7fe//��dS�by�[QQ;��n��ql���ќ��{�a�$V�����w�}���,Seܛb2m݄�3Ͱ!Ҏ�A�K���Ѝ��{36���k�]�O8d��ȍ06D]�
��!1�(J���/'��'`L<�_�Uޢ7��,����}��K��'�}��T�U�OrD�qօD�,Bߍ�)Τ5q�d������B�k�U��Z�ĕ~��ߋ�y���sX@�j�C~u������%�ѹF��:����$Z�HLI�#��!I�C�m[�Z����#�ڻ�a-�Y���ty�g��n�5�a��g��ɘ��k*y��/�h%�D�BM�����~��_�L��D�K��Y�&7�'V���K�%�]���Q���UV�MQÒs&m�R,��L�|~�C���䭈OQӐl�>)8�q��QoL9��Hi����*�3��5}�<9��ɗ�3�S0���@�*�B`6+:gQ��o�q���o��)�iLE&����h��o���8P|��j�������M(i�oP��N8*a��r Of8�k�	�%�'B����k��rLڧ#�-R�*�v��Q^��O�;���iz` q)ǋ�f$N��� 1��[?��N$S|l�)������|N�ݰ�Gs!�a`G.t�s��:U��Vڪf�]���H�J����}T���`�|��+�8=]��%уԶ���4E�ε���>����V��G��A?pI��P�n�W!8OB��5H�e��R���=�[��K+�_�3��:*��QvHL�3߽�Y�υ���"��$�	��,�
*.��Ǜ�3��8bV3��Yp��)���������6��^�G����������2�d�F�"$�Ο��UP�H���*Q' ���k���R0��_��έ����τ7�5�Ո"J����c���6in}?1ͨf6�`�]����֕-�Rz�[�v�O�r�q���л�J<�����|�b$� [�9K�2�mm39Rux]¨tw!A�1��CnBa�]�FVJB�_��f-quP����"�w�\0�n ?��Ą_~E�D΅�dJ���j��=�a�SIw�yK�#x��|@�]a���4i�#p�X0��Q CR�� -lLs����rX�f`bY���h�+�ܐ[m�L]j+�5C聾��"UfP������AA{�l���J�R�sf
���+L�e�*m'�3��W���4{O(�����W�>��	g:}�(��{���8Z�����kmߕ<Y:�5J�p����F�,�֒�:W��"�շ���!R�G�,�n�F�4ִ^�;S������@�-Szlu92�`��a��(�1��-)ux��mw�VRw�.,�7���y�uq��k�MA��x*R�k���*�V���K�>UJ��C��P�-W� ������p�f���"�c*OzZ��f�%��r`w���m�GȴÄm��1mh���ǀ�^�Kld�A��6�=*˂&���|��{3�8�}���ڗڜD��6O �!���L���r���}�OỀ�U�|��e2xz0,v��\��հc4	�
���N���^���M\-�-�J��5aD�F���]��jU��
���O�|L5*�T�p���
�$]�t��H��'0~'���S0�
��R:�Z{(��`�pJA�lx&�+��$8��P�_�S���MB�eR3
�3�	��SW	�M�)��o�ل��6��Y?�+� ����0'��'�K����*�o3�W��aާ�=��&�@Z#9�s�~"� �9y��q*H���ᢿw�ps_PS4�M�C^���zcQʓ̍���.��� ��b���@�7O`N�4��������Be�1+;őP�8�� 6��(���BWz������y"����4K��KǼ�V�5��Y+Q�����06D{?��;x:�߽�A�r�J�K ��')OކS j�x��aN�g`=��ژ�����,'��_q�믬.����}*�;򷃥��W7I��ӎ�"�JRlDA�� @�axM~�H*	���k�h� x[A+?��;[s���H����Rܘ6�,}E�ݧ�FT�bۊ��P+���w:��Ch�/��K��#zL�@&�]lsU�^�O�3a��62^oX�E��]��U'�O2j�����"!2\˱ST=�̜��֡���\ۍ~��<I6(
e	��g`�0��y̋ߞ�k��Iz,w����
<�<yZ��U��Ln��<,��i�H�|�<�:����?��.��(y>sl�01���ꆧ�k���)E��=y����W�q���O��Ƭ\�@m���HK&p|�8����� 3F4?47�U�~��ᱤ�yY''�qaS�gXn�7
�pML��� t4�=����
��^����ݭ&��4S�����ʟ��rP��^1Vkd�6�aW>U�;�	��[|{�~]Q]�PRDvX5���AG䛗�w�e����j�!V�����0�����}���)@{m6G9�}��oB�3),g�(�|P�����{R27���S������w���sGMa.�o�2.d�N��K��>�9r��~k���Q	�km��B����@��o�~�k���M�?uz`p�nr�n��̇G�d_�zot��q����A~㵮y�8"�����?W�U⫷�M�٪qYG�B��Xy�)ԅt�:� �xԿ���^Js��cD�q��}~Q��{M�@�V���`�e�q�1�&md��ٟ��p�`�;4E����@+��s�y�mk�R���QS|�#B4X�M��/e܁�a��Ȣ���}\T�fx��5�Q�T$>^)YT�i O�B�2�H}㨔]��6������/b\�ʟ"�Xg+��	''q.�_WM%�����~�&9T~u�z�w0�{q䩒����� Q����2������H�,�BK�*o�y�st�*e��L����2Z "@��;����]�����x �y�t�%l��h�	�0$`�tɞ�~�����5� ܥ>��|�!m��R�;�/���+-,s-��a^v��M��Q�8���f�����s�W}��y�d�c]�+%�@L�@��N��z��o��׾~nۊ�c��Or�����W�������<�ֳL2�hy~�6}����'�YR���q&A�����Gck��#ŸH�Ȗ�������->�߾RpU�<���A��ɳU�A�����#�>�L/��ҩmf�$��{Q���c��F��,�H*��{�ܙ���U��S�{�2;[ƇJ��1�2���qW�lu2!9Gx�.~������2����ƸX:%o�)Z�-x�cL3(�����=7��m�5i��y6E33-a�WA�Y'�w�۳�*��'�JcQ�a	�'S��Ik��:J^�9�ݙE�W2�4�3B	0� �G��B�7e�ぷI=��`���1�^9�"}}�o���3�d����������×G<��[����i��,���΄�m�U��^�}r�/����iR]�����&*����^'ً��l#�n^���I�R�ܼ$c8��:��uݸ��O@���Fc�oWd��*Js�<]>���?_��}E$��^
끅�?���Ȓ=L �V�.�G���
xV�c�3Lmt��<�L�{/�=v7��Ȩ�(����E��\����_�r���rJ~�!��84@>���R����39u	bh���...S���l��G �J5�h�W6�C=� �	f�%H4�K�	�vW�L����7���4LT�Y'|M�丘��-cj�@i��n��ô��΃�HU)~|���.�����(M���[�c
Q����C�s�4�O�2�3�"@���d�"�KQ_���h��������e��R���<��xt>>U��{��gy��?��� }�z�T���X�����֠NpqX}�8+	�l�� ���&����ݕ�+��Eэd�~���عfz�3j��r�J�ۧs$�����(�6��B��YMyJ�9�4����j}���.!�?� ��i�<UaRDK��x g,j�EK����-�i��@��[X.�B{3�� ����.����秴�/��wͦǃ� ��K=l���s�NH����
}�.���	��4������u"�?����,}ɈOD�o�uG�N~���oݵ���'�������|j|���$�٭:�����w�g������b���-i�ݓ��l~T�	7��x�qG0�W3�}Rt���' jу�*!��24_I2�Tާp������j��t��t�&:�+��f����[?%+�o|0��V��?8�6=�'sz�O ������D�T�U�L��h[ -^3[*�	i휡�X�61\h�3����h�v$v���_8�8��n_5���զ~��?�s*�p���3��� v*��E�\:��p����u&�L�
�9��}��YM��r�a���
.3��3mv�į��ݠ!}u�»��� �m\Յ1{�|����[	�@���Yy/(L�
I_�B%c�PL�H��+z-�#k�V�R�G7T=K�(JFHm��E\�sr��e [�����J��#�v	qcZ�dU�s�I��I�.2z�:���a���4]�;*�P�w�[Zc)���I����~QY�9�sE;(
��U::U]��|�!ЈS�+ �M5�"F3�I�Ҙgf��`��̀���G#�V�r����)B���p0I�J� ���I3�r�"PzV�1���{dy}�Ca���{�띐��c��ܡ��ް&�%�=�#N쨙/?�-����f�7�O/�v�ݢ}}H��Ah�'�+(�- 3���x@�kI�Q�Ӓ�[�[Ҍ�A^�>���=�}��f���PE�������c.y��P��-nNyK ��>5fT��|3���Cm�I,D��3.����m��4.��4��%Z�;��5�*b��<�bW�Q[f��1�c����'Cm#5
}K}��8�))���>~׊D��`w!���������Y����k �z��_�Bw���Rˆs���8���vf��P�}HR�S��j�����l��%.�d�����d�{҃���5�N������=�
0ZdcI�Y�T��8���A�:/��(ZtZ�#[��z�1E\W%�9ʏd�^k��+���m�%�B��*�^�c����1n^��k�.~�ᥒ�T�G�g	[��v��XGk� 4�~�ɑ�k��M�{��bCW������:��%���'�IW�#�BiZ^�@�gZ9`�u����į�'�h��ab-�A�̇��o̨PR:������z�{e���S��E�y]�Q�C�$_ =���<ﶋQ{]�������^�hn���Zs�� 	���J,��)|���d~\qIj�2��)���O����*�7����ϟ��n�E��ob\ɱ~�"���?�r�Ֆ~H�#��9x	�`ի�#և+|�%�����p���>G�{��
�
�Vc<�Mg�E�v]��Cˋ�R��;V_�N"%Pˁk4��;�^�ٵC?i�����:�.�uv�"��������f�M�`�h#�+�I�+�O�O~����\B�r_�R�'�e�M�D߷cr} ����;�ү�/��io�FŨ��e��o�+<(�bЂ�&tP�#�2��*"��EVA���/F�]�K@�6�+2u@���`v�u��J����iyr&�c���f��N��\�`�I�YȠ5��H�� j)��$KE�^����h؛T�f�+�,�	rFP��ll��T���t9��
��+�"o�X-Guy�s�*�X�u��D�H�0_�cM�𥿨R�1�.�`U�����e����[�b2'k���'6v�G�LDX3@�^Ygo�hgh�SZ1��W���^Z��W ��P6۫�"<x�j��Ԯ#�B��d:�s���|o{�����l㎣���0�UbL7����+�_yV�F� \��۲iU�G�XE�_���r_ViJ�Q֌���xI�	����^ZNկl+A�F��a)�����+c�6�l� �RFT\%��/0;}��pN��[�ٳ ��rn\2{B/��C��VP�:b�#����F^~�߲������ֿ�i����C����qr���E�fQ�},Q�8sb_��/0�H�^��p@M�����J��P��.���+���r� ���E��CNpu��L.��2B�ᒞ���.X��H��M��i�`x�����84�	RM�{����<iK��ɛƑpx�U�M��Z恐�sk�z4��s��_����;%M�v�c���;��e ��@iu�r�U��Ik�;�(�r��E��P?�
����5�lg ��b OW#]�%�|���D`I�������)��ދ�ұ�39�.�k�~7&_&@�C9C�N��@�be��C�]�d��3N�
@E�Y�x����#�E21�a��z��������w��{��|��g�h֮dQ�tt�R���n�T�co�
 �,tJ~�i��.�������zhY��ޜ��XR����zp�����G���b��?�<�Zq5�;mZ1�_3�l���y���n���#̒c������EU����`� t �z�#�6S�vg������c���UF����0e'�#?ɬ���7牊(�S�~�B$�%
7�Ղd�"^��d�ӻoi�NgT��ό7=.zG���s/>;z1��⑔!
�9����B̛�e���Fc�4�y�y� �vXQżX��P{0�9uY�Y�h�z}n˂)b�o��SB}te�W�X�\`�"v�i�X(Ix��U�Tj G,�;�@�y��$"�:�ofD���S��^P�e�ڞ1��FG����aw1]�\5�(����٢�t�
aI�R�݆j��*�@���=�����p�Ԓ3�ϝd:�5��#rk&�6|�Aی/��B�i�j| =�z�N֍"�q-��'��ټ��g�Y�u,�Q^�������R?��f��d*�"�	C ��B� ��%ޜi(��'�r,�7�ֶAK4u	
��D
��8]�� ��:�
nI�塪�(D�� vʆ���}��͘-�7�j �*��L���=���F4rc
�����S�&���ݤ7ͣ���!�%Y�����1���}�4ӌ�"�-�����|ʧ*
�A�:�|?(��T��
j',���.�i�E�JS����7T�B����c:��l=�w�y��3PBN�R� 6��4Z�11�ʮ�.����#9�+����rS-�S�i��&�S�n��2/��p4��j!���Z
ҥ>��<�8�(̓ �9���g�'#��xkIs�q���?����1���wV��i�6�j_������%���'�0��WX�2�z׋���{����LK�6��kU����i}]�C{I��D%�(e��YYl��ojm��m�oB��/�T�tї8Z`Ys}�
!t���"����9�Oe�vX���7>4�4��/�0@��9K �@�	� t�g�~�k��Q��J��p��X�k��D�e��m�O&V�_�<��q�j�p_�̪���\�����.�9��SQ��߿;�{�$��J��V��Ϲ�FrB9!k������rσڊۭ��~�rA�S����[�f,ے"�|�"N`���w�n9��[@�:Iv$�k�� �(t�3�i�/�=�.8����&�~��/���Ն����Ӧ�@��k�#���nΣ��s�s�~�탽�?�>���~��T,d�zd�Lݩ�:?����q��v|��y��N��$E]_���'�kJM��)�?R�g�n���I���d�Hg.v��./ү�=�|�´�u�MA0�I҉��lg���,$vቃ����O֞��UK�NPo�l>��sm͑k�!��^�`� 7�ͦo,Ĭ����>Ղԋ�Q@��m�W�	�̈*��;uv�W�C�|�y��Q�iY�x����	�Be�t��ަ�2G�G/�E��S;Us �փ(�P{�H&E�G'��Trm��ɸ)��s�����A����p`�Tq¡+�`i%Jk�gA��R��{��Jc�/�ͽ?xf�����(�w�}�j%���m$��u�������(>��e+�IR!w���K��?B؍ۉ�]D��O�yj�b�1-�5k�~5�k��� {S̞�������;*��K� �`^�H����- �F����5@�4:���;	�i��<�0m6:î�{'P�@;=��RЙg5��_y�BW*��C��$\��7�Pc��.���9��r ��~z��tQ�)��tb�mq$[�2��n� ��1�&)�-��+��gˠQi�g�Dw�{�ћ�3�m��5�������YM��o��E-?Թ�2%�S�+)/j��]�>`�$ds�$��sJ�T���1�✖9����:�9�u��I3��M���������\<֏4z��Mf�/�����j��W=�
�W��m��F\�si9ƙtp�8�fWv+b&����Hb�Wh*�̛�G���֧��T�F���M.�ԬC("���g�xu�BW�����N����7�빾�;��Ro�ﱩ5ҕŪӽ�2�ʰ�r�b�\(p��m�A���Rф@�6a0@��r$�sb������c���J#TG|r/W�,�I�������p�#���Q��/!J�D-���k04{S���L�c8��řPe�l�Q�ܳ>q��y�(~#n|�5�۴�B�	?�Q5�{��)���MJ��!'��{��$ 1��fo�`�u�*UD�t�j�?���sz����Q��g�Ƽ����� x��9�נ��3S9�{C��u��w"��8� 2����D�tAl�������i^�Q����G�P�e.�Vd��l���$�bB���0 $z�T�?T]��b_�;5>�eo��1��`3�.��X���S����B�" /m�� TX� o����g��g���PF	�����}���;CxMJ�9C�`|���V��B);�`�-~'��1"�?f���n�w�Ѷ�l�w����1͞V9�|]�D�ʇGa7~>/���ڵ�Dps����U��o�<�A�t�i �8i��.�8f�͟4�%���4�����Ϫ� ,=dOQ;s9��X�>��E����i���t�5��%]\y*c怵�9kwT6~�44��M��[��c��c��!p��tk�1�V7��y���*Z�_�B����)N��-,7�� <���k�ނJ���}1��ܐ@^���	7�BEP.�_P�������qJ��t����vJٕ3G�xl�)|zq�>c�����N��>�l������i��E���e�i���l�v�>;O�.��`FER<����$��j���W��5=n�����^��q��ͬ�/5�^˖�.��ߌ�m����Ϡ`c�n<:PqE��|��`=n�x�� k�a�㧥yz�ua�hym�&A5��o�9��0���n�y�R㙏7�|{^ A�iG'�Z�w�]�(:5oISX�i_|��o'r%�%�?�7���1z��/.�,��4�Z��n�c+�V"O��]��y���8��F��j��e�X�$o�Kކ��;	oFZ�?k~ �|Ac㞴o\ҍ�� �}�N~�^�32��L{ �&��[��g�*=��{�,r��]_�j�M�D/$�\�YrtY�TÔ��r�*,�啔#{�w��G�=AqrP��h[�28S��]v�]\��.T{���zӹ�Pv����{li�pT{����j-��%��p*��R�X�� s��I����ڧ wM'�0�����P�G�N���b�i~J�{92e9ӏm�:��Vj�#A�2��C�\���Iw�'��dV�u�=Y��w7�`�H���[�H���ܵwi���PQ�y�C�V��)a)�[��|��µ<�?x���r2؞��+a�>��� �j:Y��:��8�/ɓ����^ ��,�o�4lEgU-CC���o�OP�*V�P!=S��2�/-{Y�F�?&�a��ˑ�Z!c\z+X�U ,����:����|�/��R6]��nJ��p��]Tl�����T#f컔�d,w!P��'��t/��O����׼$C��(ԇ֕!NA5�"6J�֒�8cb�@O�7�^����Ts��zR9�R�mB�.:|>+K[�v���2�A�c�~���	��r|����O����=��l>P-�vV�P�±)���x]'���nVv�'��������{�d��R�<�b�}�%;�#`�ܤM��ω�c}�~�#��������6��F��ږ!А���������2?��yb����OXW`M��H6e��q��<�\�L��Y���?��Z��k���W��` �Uv�d!�aZ�r�9�W��������W=�c���@t1���R[����+��L�	�:l	�fH��՟�I���|O�%��!O(U��X�����$O��}Sh����#Z�U(�i��b�m���༳�l��SFS�E��$Sz�h]�F �Taz�����8(q�ܮ�ߒ�Wc�К͓�T��}�[*C�۪���bAh�18�����R-��Fq�!ߎ�ϰ���K)e���`Ǭ������I�5�w�.VД"�ībmܖ0�%��t\Z5�m'�wqP�$�o��s��8�\��!3~���q�nA�M q*���w�,���K�<_�>��Џ����3��_#S7���(6�CluiW�Q�Ak�e��ݏFI�E���j�i��ꅊa;G@2
�� ������`\`u 6�o.�m��T<pvl�f��{����|�X������rXɈ!+��SoI��n���vHh��a�>S�x�e�3D.��/oJ$6l{_�dl��UB�J��X���KB�q�(�l%�v�h�O��̶��G<a��#5J�P�������|�����_��;�3�5�w� '�?@J����V��y�"&�(eBۺ����-���K).��0m����r��{�>y���8s?r��=���
�Π��k�Uy��Z�a��6P<��n���U4��R#	�P;[6߄yN{`���T����f��cP	l���
P���4�Ք�3����y�T?���Q���U��M�LptoP�?0��W���&2�_��}�T�<�>7�����Ri\�2�;�'��a�_�f�L{�`��� ��xՃM�8��h]�F����F��MS���<���.�g<�֪��L-�]� X.X����W��"��Ji�<Hͫ���ϗ�!>P*KP��|���X��R4p��f�n�J������X��P['���V���v��=:�����DfP�����9��[�K�����.>t�1���ꨪp�"��ު�#Yğp"<��?
��%��~J���9�&����Q�dF�>�h����3��i"'0�� ���Q�v42l	=��D�f�,}q~ŏSKl��"u��!^���`Ҵ���&ur���+1��'�:t���D��,�>� B,>�O;E��f�"������d^��9i��26CG.݀#�[f�$��MG�=�T.�R4�
i~:DÈ3?)y=�}�[*�M!IC8d�q
�W�Q�����@hr����)e�t*0�&?�>��g��̳So�:��q�+�I��C��g��
K-�ƪ�:�5dS�_#wD������]�30yF҅�5;$�H�o�O]�l��������a����{, �y��\��T�k�l�HV�%K��:���@+z�{$| �;bm��-�����%`^:�)"�Vf��ԣ�~O���I�)h���;��ڛ#֮,�� �M&�$a�x����2���{"�����ә�db;N��ϖn���Qh�ӊ��ep������[2,�F� ��w��lz���ig��>�\Ѓּ�C�#���1�ձN�Q�r*��kW%� �*���R����	;ؿx���c�Ύ}Vo�����Sf�b̃��L.[���"42]F뇪:�}R�ٖ�>o�Y�zk��T>Ks<w�L7�+��Zy��h��6��'�Ws@S��Jh�ב/p������*w��<b����܎�8�ȓׂH�9�`X��Ha�&�M+��p/�<&�2X���]�܈��/���㲉�&��`2��L<��8T��BRN���L�^�R,H�$2�n8�\����P��yu�k�T���DO�G�>~N>|{K���U^ �Y��
����F�'ꬭ�7FI�}�]����,�߻DǄ,�� ��3��nG��������m��(Z�(>e"��ƅ���	;�Y�Waq���͋	���U�yg-ήX�]�A<ϲȲ�L��c�c���v1\3���
������"�U�;�R����v��Ժ֫�S�<sN����c�>�1qp���h^q/|A�5���yzT\|���eg�d=N�Z�Ɲ�R��Łm�݆R�A�qa��O;�!M�.a��B/P2U�'F-��y`����� �Ez�s�->3���꬗kr�Z.[£�a>B�8P�_r�l�sO���pYT:���q���N4��Ƿsd6��~�31}�Va�V�<Zh8i�N��i;ִ��ld�S�R����R�
e�0�۝ͱ���S�boE���21J!�}�e�@��_������	���Է���B���D_� h��)��1��¯"b��O9j�l �jm�Ƙ.���/s&/!n�p[��Bgz�|�W�Z��6c8�1\x��-M�t5�b���v�C�iF������.��*aq��I8���N��Py]܉"�0�|��.)�B���[����UK��ꤱ�-��F�I�F�t�pon��k�[y����9W��F�˂�$1k�'��4�_�Ջ:�X��4�z�V�6@���eG�������������TD�~�lڎ�*�w�����TB�'ZV�@�g�mH��k�c� * ^U<bZ* kJOG���q���~^�n�$5<r��g3�KҍJ���ڭ�N���~��݀�z]$�/��#���~����$�tL)o�(���տ�6Ţ�]��e=qK���3I�8	C"ߏD��Oe��Z�8Q�i̵ ۝i����>4K��+4HKO'3��X��?,:�b��	��bA�-����|H[g���zŋ�3�c�H(��Q�;��᫶����G�5�ˢw%^�eҢ�jv�nFD.FLw�j�OM�A�zKex���Ǹ�ˉ�	_8{I��]��X��#]&�$����.�绤�> �%���T��-�W�ɨ����~��ޕVn�7y�V��ђ��q�H{L�Űn������՘�&M4���ҫ�#�ñσPeĘz͕�#���ð�Кf}���:D�HOg���%W�$�5%=��g�)�%~EG�>֗i�<��5Wk4؄��e�)&�Y�Dw=f�����g����#���x6��g࿢}����%۞�G�!��N���GӚ�DB���I�aO]�F�L�t�1�:fM�:�|ι��Rm�����;W�bWj"M�6�Bmg�A�3��D�"�Ov"6���Z�����4���;&~�$6��8�:�b�g��i��=>���X���4�R����&_-J�9����]��^Q��!��2�D]�^�K1>Ŭ*{����bJ�R7��a�߼�sr����m��W��I]�;��a��kE�82\������j�c��+q����[�ԵV_��b97�������g�5"��ޅ�*�`dPĽ��;���M��CL���4Vr�/��c-�d�δ����C���M����]�n��wp���8�6e�lS���}ƅ�p�jJ	�;�z���~�t�AG	!Qp�3~����i�紡p�X�
��a��G����6Iq�m��f"8h���%0l��w�N4^j��nCY�-0�Ƴ���R��(����[�r5C����t6fV6�6UаN�=�!$Z�	���5M{.ֳ�W�R(32�J��o���r��h8�:1�J�N�N�b.�y%��>N����﯑��r]�p<� �lnY#Ӫ!�+�qY��p'���b8}���^��'�=�~��������'rѯ��/ٱ�jO�5��߈ҍ�ӓ�2�G5�o?�P�.yP�V���jޤV�bUtѴu1���s�*W0g%��E��3��!�W�F��#b��U�y��%I�	ʠ˫;g�o�'k6Ջ|�a%�|r������8��~h��La�Q/d���<����=��Z�ܭ0���^f�V/��*�`����Pb�z	��k=�GZz��\G� )d/U�r�Կ-�s����Z�K7zA���}�)� 	R��$1{�1&�S��w�2�¥���I��j�T�{N�nq�\s��l�T���\+q��0��/$O�<�H6U����|0�4ȓ(2+#�7�`
:r	?��e��Mxss�C?���H����8`c���{�.�d~���/��2��/����h���+��#�T=��,!����K���[Rm�����[�"\ _�ֽxR�l+
B��6� �"��"�4���s���$$T����l�3�5�{��=M5.�U�v\���❭$�;���ݚ��a��H�~�\h)�C{U!±�?]��1��,�n��X���ښTP8TW�%���.pQƎGZ�S�N�x��?�F�
u���2����h�����Y�LSr�	��0, ��n���q��ü�Z;�B_�ԃh��N�V~rȁt,;�({Y�����U+�:gV�϶Q�Il�=�Gۯ�[�]K2�@ fQZW��C���oTP���
�-��d[F��{�k��`9�����/)�y�1��"�m�Ah�
�F{�a�XZ~�;iG0�X]w�o����0hA�*�k��_%�TW�+�<�%�?6F�m�]N���g��f�9���bNĲ��Tׯ�Xw棯��S��)P�;QѦf:$N893�6���ћ���ӑ2z��}�?|-�y�Y�&`D��zq$o�ܵ�#q��od躯�]쓦{��#Dtga��6`z�����ϴ�R��ts Yu*�CP�6x��Vs��ؐYKW�:ɭA����Y^%���=�O��э.����|\!ld�Cږ���d0��}��E�\u!�[�y5����_\�e��g��g�-�s^c@�=���c�k��b�Z{KO���Ԕ�]��eX��
�{����
Q:�	��ͤ��x�낃}h+A�}�v��'S�IJ�{�,� uu�;4\qꕲz�����l����B�%�7��~N�g�z�����^���x�����<PU���9�1�%���k,<����o��bQ�S��A2P4��ͺI�4h���G0qu�Z+s���Dd�r���A�(��~�!��u�_��f��:���xt��R�_֭Ȃ�5ڛ��̂��I��uc�����g�Q���E�����)Be��_�3I�q5^���m�q3LAԍ�z��0�9�s�F�*��$��E8	���{��q�<#�$}n�v[�#"#g�(�wLS[���r+�Qv`���E3�W,�w釾$h�܆7y������=-�o�栐��V(z�)�����l��� 2�n��Wx���@��ɉ�A�
ߘQ��"��Ʉ̻�� C�kԐQ����R�e�>�ǒk�Qq ��!�/i�}﭂a��_�W�jK����X(�9��B�3i|_=�[�p4���+��o���>w���C3�p+%�W�@r>�� ���-EKֺSY̛�~��ȝZ��� Ɍ蝂EBf+��#�ޯUw����5��c��TI�?��l�����\j��W,��1�| n��1�(+�-h�Ǯľ��:B-X��v	�����R*���xE eu/8>��מ6��O�!�"�2��X�B���E��Ld校��my`D#i�k��B��"�V��(wޕ{��Yн�1M�^�8�V������"�?�k���\ȉ�	j��`��-~�Q"�A��{R���G|kCv9��'�KH)8��]�a�����k�`F�m@ʲ8�c�����'(�)$_x7y4�^�0DQ�>��ZrG��tZ�h}�|:2�*g�n�!�RXa���eR?���9�{����Q] �0��{6��[ =C'~�����[Y�]�c/����[Q�@ݭ���#�k}.�����e�Ć���ӨI�z��S�&�����Xk�����	i�I���;J:���<�"����I",b�� x�r�}=����u�r�j��'�nz�"�dCp��_�w�љ����j�j->��יN�
/�N��}!�Ał�Z�1?O�\Z3��{��&ɗe�lv{� �<�;Hw_�|.uVָ����.Z�u8|<c��5�Q.��:㳲�L��鵞�9�eP9���US��N9N�e�Jh�k\��&�Ǆ٧&�8�D@݆�OQ�+�%&*'�MF��*���w�(��4�>�~vgT�)�Iy�Xsy��}�����i�)���0�W�!��%s��) �}��&ǰ��0��K�<a�|eL+J5EM�dX���`[����r�U�N�3LgsZ!���k������4��S��Z�B)�(���bvGxb(��#�Qz�># �ͥN����F���]�{�lD}F~���EI��� ꝋ�?Ǚ7��)�m
�v�+�W�X$�,"D���Ң�h�Z
�{W�W��-�.w����4gX�ΞmL�j�����:���2���&�<R�]�"܊<�7�%.�<�'��i��e#ʲU�����>����-�ܢ�^�bxf��K�Ŵ�E19�5BxgC���0�αK�	!�*,�.���~��@�P�SE�5�� -�T�� �,�) �������wT,��od8�f�i�O�nEW�����k�o��� �u�3�ꑰ��E9?��3�����z��]0� ����^��V�������*q��$䅋꽭w�u�K��wW� 	 _�����i����eUQ��͸|��yfp����<;Z����{�	g�1��B��r��إ�!���}�K[�1�d$,�J}O�vB�Hv�$�/T�N&\�1�U�#^�I��,}V�r���^$�p�*�o�W�ޭ�4�/t�=1S��:G��T�s���nS���]S�	x�ӏY{F��XG��s��b����*<$bT��7?�ȑ@Bt����z�3��.�Q�n0R��Kx$t
���P���[��a/�X�T0�X���@T
e����E�������\���j���#��(s��sKa�?���/���I��G�����>K��7ky?}�"�+�R,�*ӎ����̐�ij�{�KZS�����i�ZT��$��$�W}�\��D/�9��W?�9��aE�=���T��a�@/�8ev��U4�l/b3k�D`�79�Ғ��+xA�An�R"� �}�a�,�Ȑ(UZ=aI�dp{�Ѿ�d�N��84�FY�jrK��K{�>E�����O =ҷؾ^?���U�GV��s�ِ�G�@�1�xEO�$�]`Q���hR���z��ń?�@�t�1���2�v�:�8g~|�V���p<0���D����B��v�5��s�e�h+o�#��L��H��!@]���|����I������E�G��7�H�n�y;�k`�4�R�!�e��:d�O'<)�r�BE�l}{�C��y��5�9�٦��SB�s��WG;�Te�����uO+��$�g�H7���4���Q��i��8��O��95_��h�)�I��{����xϙaz�^@3�um"�m�g������R!%)�l�v,�t=�ǔ��f�Jrd���R"������D�z��0����D�-L��'�����TM�x��`���e�$���'D�x�CVT��Q")k��+-VCz�5�ӥ��A=-*�zP� Kl��p�4�6�cv1��ݜ(Ut�_�� ��t��R����o	�؇JM���I�-�R��o+��{8
�R4��qc%�W9v@7�4��m#�ǧ��<��\��1#a��F&-�R��jP�u�3L�E���%<U���߈p�CA]����ESx�>�_�2��� �螊�GZ�,c$�-XI{H�T�J��@2�#iM,G��A��0~��,�p�-�����>zm/�
�=�ȏ� 7�FP�XuO��g�%��QT����f��9!���A��"-U"t�6��c�_��v"���$RZ"۳S��RR��ny;l��-^�!$�yE�9o	U��Yr
�S�[���1�Yi���a�l}=��H�P����.�2��}�>R�����k�t�BQ�7������ӊӬ{@����P�-��ڰIr��H�TΝ@t�����_Y"�����aڪs{����	o{Uc��;���峸p�NK#$J��A[T�3�L���O�ʋ��oLY��;��C���Ǐ$��N��If���q�A3}4��B��{ H�X�X%[pS"pj��fmW��c�/�c�j�V;{�̉n���������q�4 hi��?ĲC.�1�=2kc	r��@ڍGTh��� G(e��ЯR�i��r5.������E��EkO�ղ�pԶK��I�b�\�uf�3$Vd'����@X\!��W8l)�-�����@�Hbڻ�UB��6Ff�h�
*'j�qzM�M�z��w��&F��N:�i�)��I���1*7N���I���%���G����;��]����0e*=��0������DS�[��:�>'�:�l��9Q��I��/�Z'��^,�ȑ���$��ǥ�����F5ҖTiX0�X�vQ���=)q~��M3J٥W�Z�m���<��Y��Q�h"o�1ܬrbgHm�����\,s���킇���٢A�g �j�a�M��^��=���d�`�,7��%��~�����2�zI]'�D��¢ks*"�9�tͦ�qM��
?������P�'�$������b�D?G�Iz��!Q[�R��f�Z���d�v��HK��A�v��;p9��B��m��heH� 9ѾÆs��w�/?��<: �]8i�<y��M�V�����Qnz�UW���n쐢��ll�/B��4�c?hh	�>�5C�}�d1��ZZ�p�âl�V���!D����jU�fH�Q%�Ӄ���`�g�����Xv�d�1[chUO3�#�<�S�u��e��c�`l:�a@�+�Rhs+�hܪB�3��X5F�>-օ,����i����[�<>���_��b�݅���]�!�}iA�Z�j�׮���e�\��d@���������UXI��|�5�Cea��L�>�#����P1
�#T���O�V[�*�FF��4{Ҫ�z��1@��%��EyY?t(��h���Qy����a��>����0ճ�^��Q���I���}ԧE���`�S�U_�2�����^�~���!���5.�\�Os5Bi���<���B4y��j���V�e���J���T�Ϥ�nז��aqY0)ֽ���j�A�ܯ^{1A�B^�%�d������F"銪\6	�vk	_����&�..t����*��Z�	0��l��{�^�aC؄~[�����Ub6�C�>Sy�`A1�X!�୲�<���'H�燴z���r�0��C^k�iJ8LԬˊ[~������||�MW����/�U�Yf1aQ@'$
���9��-�jƂ��7~�.|`��{�6�K8���Y%sf�.�a�����@�2��.2j��'������蝚���*��8���fd�۬v"�c*���v����q��x�>/ ���w�[S�7|�rf9���rc�iR�C,_�M�]8K���{^�Sru��536I�BV��8%Q�<WLW�$�&/LV"�F�r' ��4T�hy�g*�����{ �O7�S��B߆\�	��W�t��]�t+���h�i��<v�+Z�e\I�;�8\ڽ��L��G�<#�T�����}�ݧS�u��+~���׽c��/';7�I�����^ڐ;W��_��Lm�o��۷}m��]�j��ꀢ"{���O�V���Y�8.�Ǚ%����)��ې�p2����G��E4����&ĺ�����n���t���*����}��=���Bp�;��m��n�Z�8 j��v����]�{�_)L�`i;���eH��Dx��+���k攱��b�-&̘R��p�X����ՄgBgS�^�|=�N�S�uZ��9��E�F��	շ��������U2���h}�_U/<���~�wn2o/��֌U�n/�kJ�@f!�<3�}�M�_"��@��f�b�V�/�@ۿ�$s	���xT�L<��[}S�i��YO]������1�V[>�j��� Ys$�5�D��q�k �7���S��t�	�$#��Z��4	L����}��T������@>5�������!�sԜIq���O.{�:B�J�k�4���j��_�ubd�Hl��8D����'��&/I,O
��*��[���Nt��ȳ���=@�pu�	 ���>󈶔��S��+,|*��hOY6�{���s|�+�q���V�-y����T35<�W��G�b/=&��/in$V��y�ėS:7�,���Q{^�_y����]7aR<:/���/1ib��!��A�h���n4J��{I���q�i X�k'mg��;�D3�A��N~iƮ[k�w�0�*��m��h
�'���'��>
x��U��y���Z`�.��u�a~&PEt�����.'����Eu �����q��M)�|%E�n�ծv���˖	������\أ�>7�&4��b>z���� ��ޣ�Vk����W�!���-F��;�eh}������~xSҵ���&±�%ʯ��ږ���L˸��Z��Ε]2�4a-���4�|n9ݦ�D7��,���Ҷm�8��Wy�������c�PY���;�N�p���(�/� ����oeq<�	>�F�\y�=.q�@�ßz�7ݯ��1�{��H��}ոX�'L�υL�Dl!�c~��~zH�,��k��֚�S�3z�C�� "��A��)g�(�2�m"���9&(�ě%�� k�^
!�k�a�'��+>�tB������}'��ѓ�S�.�e3�7�l8ɬ�Q��[-ߍMuC���{>����,-��o,���*t�z�����2�SZ�y�u8��U!�qa�� �V�p�k��,�����ca�Mw�S�����l*㊊�|Q)@;5DB͊�yc_�۸q��q�x��iW���>�T}����ުQR޳���,���"�O�5�&V��g�v�-
��=��c����<C	O��@�v����nh>a$ ��#���a�@���w�+F��=��!����LJ6�I�;�	 �	�G�'s�>U	rSQY��й�^�ި�͐�;״����~e��I@����f��.I������y?�I�(�Wq�qe���9�*�7�*�Z�-��'E�M��+�<$&~�n N�,H���Q�S�>�=D�v炬1��k����)����,�NL�;�a� 
oU\�T�{��`'"�3qp�y��SI�)NW 3�	)r�B�K�$��j�7{9���s���$���uŻd��������|���i���'o��Q�t��[7���H�0�`8�@ĺ��i����w|���.#�q�B,t����.�qC�κB*3���T���7�[�١��W�������d��oq�P�ry+O3�Q1������`����DNc��?ҩ�g٭��8M3��k:�ݍ��;����9."�*��Fjd�㨓Cm��)
hL�t�N��H%��z=K�x��g�!EW�LWevQ��A@�U�h� W�������i���x�]d�Y�my@�.��ֱq��_S� Xb��}��޿�<; 3�B,t�`w�A�1�I�a������m�/�-� ,Q�jJ�ѲD����]���\[M��W�7��eiqyy���D�P�Ģ"?���0<�K9Y���C�B��B芽��={L����O�W缊d�>V��B��+�3_�@U�B����J2b.��ï�U�G��X"}l�y��7���=j��Y��9ڈ�
Ϲ�׋���_D��jg�޼x����k�yN+ȸ$���x��ty0�g�����+S��7	�u�U��sODaOK�:��L4��TKwg]�܏D�R�qlX�9dG��WR҇��L�����ܻ~�s����9i�#���������G�.�u�����me���;��1 j�S��N���Af��wL�\��$q���Ըܰ����Yv(0e�]��ג�	gŘ  ��jkCX!�d^B��|�����tW.��W�L%@0�,v:`��y�A~��)�"�OQ7�jC�����h�{���Y�;}��ž�{��l�G��i6h@�Ue�㫸5��E_���ΠATRX���-榜��1[��v���.���_�q��s
������H��p��E�4z?�H��9+*GEڑ}�A"�)	(a�Q~/L�� MBZ�?���UƳ���ƙ��蝂'�GY\��^��/�-VW�U:-�U�l�ا#]�赀����P8"�w �2q���`�̡,�.��SZ�!�(A0`�3�2�7�;m�@��0��f<{���ͫ�R�򔷘9{�>B؛��	�b �6zMd��xׇ�Cz.����R��k��̜��	�����>!��#��S�<��A�ק��S8i�XN��dT�����EJO���?\R]�J��6��~�u�?��X?�W�.��r���zz��@	ʪ�nnܙh���5Pzǐ�aV���~/��&�i�k���je���DL�=�RW+]��D7`����ᱝ�@@���E��)�+���R<h��H�cE�9�\0��W$�ܺ���L�MP<Sp9�S���S(���8~C�����ĸ(���� ;��'�'�%��&W�K$-�0�[D?����ti��_�쳌��j�e°�p%KT\����|�����m��byrp+�h�z� ���d"�[ �����Z/G`�G�3�u��Y\�hss�r4��(�LyR���%����O���/�Qf�DDO���h	h+�*�~��v�)S{g�.�B���[RP�FL�j4�3Ơ6��ʰ�m�ȅ���݀�u�Y �J0��`�0z�T9�Ij=&�V��RϯǉuXl��ԥ�
C�u�`��
�]�2FKbR9���	U���i�r�kF��y�Ja��4*_*S�xwHl���m��n��	�-���)�N0�\��_���|{v!�N1}a=�>�����Z���C/fh'�1��%���b�_�}�ڢ�c�j�	�}S`�{{���c�[�������c��dz��	J@�+
,�'p3vg�g�����a���
�)�F�7���~e����%Ɔi�?1�U,�3Z�#Z/��}��^�`�pH-�%���)LٔQ:��\�ᇨR��Ay���� �����hqD1HG���M��bz���#`?|!�m��]��L�p�3Mù�CĽ?�p
bx��?4W~&�A�� �n���
>!&v�S�`�y^b������seB��.�%|
��N����gE�ʾ.����� ���k��Pj��?� LI=P����G�^��Suz��q:��(��r�L?@z���JjU��a��������x��Pl.���ԏ���{t�߾���n��3mY "�F��RoA���z�|�(>�b�_�U�f�:�%�d�6��~)P��+�W뻐Z>�Ʌ)���8^?ۓ]o��N�w�X$i)��F��N�L
��)H����I�����)I���5$�,7�,���{��=�F.��քə�����zN�G2��Uo�#�y�{BiJB���]c�����9���V5�=X��B
����1�
��y{(A@�ⷊ�8�U��nJ�}�Fq �a�mDbou��06��x:�z	-:��6f}r~����vU�oBa���t5iL��ȬXQ�zlP�ɰC��0ǆ�̑w��^���%������Nc�]�5�^�4ǵ��-�����AHF��`}סtE��d��2��b��%C]g�������YZ=�`�߷�K�N���0���A
&���F��V6�D�+���ݖ�	�vG0����}@�.M/QCc�o�ɓ���[�?���U��h{Q�{͍u����C/f���_Y��D��zI~���aQZ_��昰Y��?tt�¡�3����b�׌J*VUu���-�,k��R��*�qL�j�
�\��}��#r��T���ܹYF��0m0)��F�V����_�.ӜB�E�����^�h��@ڃR�8���!%�v�[1_R�}\���@X��xkߏ�6g(�z�v��5V�P�0���5@��j���B*��h��e\Y���%�y�ˠ��c~"���0T�8�?��09
�ጮ��b��Bpm�?a[�xH�i�A�i�9�(J���V�_����dt<��
��c�'��|�0)t<;�f��Pٹ�:I]i�A��y�^"�u��9�3Z�W"�r:GE~է5/-<d"�N�īGb2���c}�isD�"�m�)p>� ���~���kA�n.h�;�#y�rlU�3|dڅ��t���%�Td�H#YY����sȦ�5��ۋ��O��Ɔt�Eޱ�	�D�T;T����Yktn�/��7Ѣ�ިf=��'��#���ZtlhB������~�&�����6Nֵu�S��(�=�!��TSF��;�Gb�](S����硷ˑJ=��ޘ-ː,+�m^�
������),\w=��;���Ya��"�m�/�@5yJ��E�l�������i���\�dP�|���/�1C{�C4�
�D��^��kQ�W��?��O�t*��$ֹ��9e����[���N$���NNXks1�-$/���B��Y��>s���d�^��
����y{���I�O��{5��b5���m��G\�#"���f�>��Ĳ-��C��c���k���Y�J�v�(��
$6����&V��a�Ӗ�pq6P-��ۖ>�xB����0��0B��W~O�/����!3��͛�M/i[v"R��sH@�'��^�=������w��/о�rw� .��f�&m3 |j6t�x,�}2�	i�"��/��
y03����9�y.u���JA>H+�ѓ�G��Zɣ�uα����=�A�b��LlM3��lʧw4�"X'Z�S�r��*����ٱ(B^<��m�HW���\���k֞?*�;�;��i�O!\��;w�g(�$ �OR�.V�3]��S���3\��Cs��/3Y���fY{��f{�������m��
�Ľ�܂�q�{�q������}�4ښ��Z2X��������GYr_aHsY��q28:M�H7���N�(���F�"y9�ϗ��2I��]�w��c�\�R���a�>m�Sx�\[�w�&K>۠;�!��cR�"&5[�7|���	��`�M 2�o�1S�F>�@>Zo�f��ԫ<B���������$���H\@5\=�����tF��_�F���/n�Qxj2����(�N�N����?��t*!Ǭڐ����Sw.�}���)�NV�9���uG� H��3�]1��uj�o��x@j��L����v?��as�^b6��sk���y)f�k�T�u귶��;�S^s&��eZHјJ=�W��?��*���~���QN��Zn�9u" �,��.��(��-�¼:�7KU�nK�h����*��lE����6�Z�������f�'ge�D�	`KԶ��	$�����(�z�*+��b��� �Xiⱟ�DX?y<4h��]zҳًm���چF�1�C;���������!�j>Y�������o����~@�̟c'vBd{��\�9&��QHΛ�;o��6�n�֓�z�uG����zO�N��w����c^h}�ԙn��Ul�Xw��II���bx7�e��w���uq�D�\����P���{�#��}%���^P��sm��Ξ:D��Z� �M����߄B����7��#[*�B�8�:4�E����lXx�����L&��GR\l0��X�vY7'\\��=�oo���v��۫�;E��83;=U��5-Fz=��<�Y�ʽ���K�:��<p�w�@��3�0��7��x����Q�Y��%�ʍ`�ņdܿ�?���P����!PV�D�H�� �>
ĪS���z�I�z���OMi�r�A&�3�@�ɠ=%A1�lqm7�nI��!8�ĝ.9ш/�ͻ#����j�٤Hy������������'G��.(EC_!���y`3�@�Ӷ������0��,��ze���w�X:'�k�*���ΎJLX��`�0�4r�w��Iݓ`����x�`����`J���M@�0�ы9o|4��r.�@��B��?vI�+��s+-BG�\&Q��=//N�vnD��?�q����ɖȢ�����63�����*��!�K�i��[#\���!z�L#� �	KD�_N`Lfºp���UWU�}o#��U�d��k�}�GܾSF&r�o�f4z��a�� �6��TX<|1���)"��M�Q�Ȃ��EhęH`1�^2���U�̻����륳����+��÷��۠9Սs�˹'ͻt��uϐ�����]gv��^4O�/d�,���e�Aj�q���A�,�9�EmD�Jv�L��NK��"�
�D���?!ٝ]I�� � �c���vb^�l%c�i=�J���%Z�ǀ02��Me�)�����/��|s�N}�VN�Pg�;_+��-\�Ɯ�����|4�5�C���w�����r�t�ü�-Xl>��Io��=B�\i���ĿP8�f��@m�?�g0g}�#�n #<$	z,ֆ{�"��h�8N�n����gu���h��|�X!����L��X|c���,kᆈ\W\s�s씚YB��Cϰ��x����/��G2Q�1L	6o:-���w�:�5�Iϰ~���E��Z�����>��F��,4�(��
��:��*��߀�fHW�[JK-�"���i҄s��qi5L���r��{��$�0����e����'�r��L�.p��b�yG�f�V�?s���XUjA��	�>&�qf�j���Ŀ�%�c�/E���n[$��hǬ�����O̓��Ea��N��m���$P��3)o�O1]O��K
.׀(���b+�wuR��	]P8B�&�OQ$�=��i}Z,��	1u�F�<U'V����9J����/n�����F\��lk���D�xxl�'�]jց@�Mqv�Ex�	�4��ͥB�9��i�e�-bж�ĎN�y��*��Oe{(�BN���K
���^C�vD�w(�;���Kp��Ȋ�n1G��џ4�����%�i�-S�<��T��^�,m7zE;xZ���)�|��@(�kg�б����Y�.�`�����(�%]�7�Υ>�;&�}}3΅���+�ÁT��wS����ȋ$�'��j�� ��)��͌��`.I}���(7ܲ��Gl'���~���ft�m��ga�m���{� 6�g�����ʺ�Z�:<a�i��l��@���hf>�|��ߝ�E���}�nϋp$q��2�`/V~�����za�D�!#�1t��Q=�[iY���飺��ul6���KMY�, ��' ̇�ދK��;�����n��8�� ��� ��M9������|���6����V^"�=�Ȍe`�?��lѰ�e��T��M����T��k��yZƀ@�3/�����u^R�l��-�>t�\�����D^�6եJ�P�z~G "�2����vG �I((���5Q\�llj2�ےIH�D��R�	̛�����I(�bvy��z{�ܴi�6"��+U6n�q��v|@�ޫ_��Q	N�unJy�vx�L��/�kr��D_Q��:��s����B��L��8t1E�@<�5��F�Uvo�?ej3ݙ�K�܊)�f��uV�J��>�<�.Äw�i�T��f-ӝ܇3'�^�Ѥ� �=��k���@[��l���p�/�p�|�/��b�7ը�rQlS҅�6K?24P.�,����ĢR�%=�Uh���\y��>1�h���:ZR���=B�,�i��J!�;��a��n*N�D���n����@�.���C�C�՜��<
)������� ]�?��q��N"����?�Y�ؐ��rP-�����~W���"�7�$	�xQ�#U�]��V����E�.���52����� ���YҠ��.�	�E�A�k�b�u�ۀ_[���y%����	�%�u�v�
w�4��*v����!��8���=�j?�֛W���KD�6���]]K����i�pȭ�J� 	<m~�޸G�ԆM�t)����_��
slBX��ݢt�  ̉n !E�w/˲�X�D6.QT��v���Yz�kvI1�r������)� �V�0��a+�G�=2JC��%�{��5��	O����-���<��x
��EU�a� �)���j�q�{cN4(,�G�O
��8A��F53�1tw�p,�*�jCF@���5V�o-�p����RaVܲ1eXRlc�h�ͱa|-nu���]#a�K�w�Ca�Ⱦ��d\�N#k>��_X��X���B3AΨ����j�/�ɖ�4$�J�R�N}ŀd��Za7|�3�Iw��Q��7���3ff���`�k~*�G6D24�+��A��9Pp�ݶ�LC��Of5�����I��� q^_V�z@&��3����1�]悩���T��j��w6�dUp�aA���@Bf�����2~�PZ��ȊI3щl(�C]�k�g5�zB�����"�ၝ?���c���q�F����*P���]��c�1�|@�kt�f,d{�V�<a�okJ+ ��3�m���m��R��s�6��ʂ�y#���Q:�Y��J]X��(�����m��1��z�gJ���茰b�*�^���gl�%�F*���Q'Kq�8��g�!(��5�������e0M¦�v�2�����Z+A}k-�j4�
n؝�$n1���73O�8m��/���f:y���GgՕ� P��Q�"�/��,*�Ax�-�~������y}�
�#&���Q��$����b��X�z�ҩ��L1�<�>v�a?�+��.���ttR�&�c[W�{�^`�Uǆ�wdj������B�FC�9��$�\�@��#�D���+����:��I��5t�:gʿ��ئN(k5ZB'�ik#W}3�R?�͓���.�o��8�� �T�yv�dMv~��go?fQ+����5|���Mv/��h,�mG�v�hDH��R6���:�V�i��N���0|]���sJ ��^Ic�ς~�3ͱF�ϊ�; lFA���y@�[hH�Z�:S]BǌJE3�9;����8!����o� �����]�6� �j�p��|Z�fDh{u68�QM�'I��^��T3��HM�x6�z;���%)_Bn�������ZR"ؘ�z�}y�a�D�jxMs�x_���S�)�Mug�T���dhu�}In�S#G��@�2�`�U
�Y�ݍ����o��ڮ=aP�����M��С��0�t�&  X��yJ�MN���6m��/�)_��������:���i�AiCu�ϲ$�
Ah xiR��Q-�)5h*}"��	T�3Xa��U����Y�y�V��fq�ː��&7u7���̻�8���a�<}H�1�rw_y�c�3,�LJ��p�!s p&uP�Pf7A�s1ux#2�P�UV1���v�#�#�*">��]�l��P�Su��'��l5���hv���A��g:3V0�aD���tm����8n�YxGV�e�ܳms��9�Z���e��ŀ������Mh� �?��((| �۞؁�s�k��R|Q$���Ƈm�x'��*���@̐���K�����߆�q��r�	j#1�%�E�!�h<��@9Q��/�\��V�"���^�U.��[N��c:�G��i��z�>%�O��"t����""7(�I,6RB��A�2\���ݤ���]��-�YѸ<�?q�]d���=��a�L��>��u�K��-!g�A�p�aN�C%g��V����4�I0���o���Һ�����I��1�kw���C&�㝅V%�D%X�yZ�\��耊�1}�Q�����僳3��S_��2��NH�]��t�������i"�y�X�q�K�EX��A��r��d;�Nm����+ϗ�∦�w.�?����Z!���e�%X�����WZ�n��$�}/k�_u��R����E�m�K��琬s��}�"�=o�U<MV)��7�ѱ��٦TV{7��ex|�oM��~yT<Ӯv]��5t�Js�g���H�k��w�a����
|�a�/D��U{F֘���7?����/n�Ĳ�E����f����!_}��dԊ���� Y��C?E� � M���{�Ą����/	c�͕������uM��SFe����ك�&�ޮ������7<�H�,]1�ף�خdन�Yj��d	@M�G
�5x�Y!��0�|�������@&b���/���ZW�2Z�rQ XIɛ�2Wj�9�Y������I6�Pc̞y��zJ<�u�T9�+��|಼82L�,�	a�M6L��<�P~�u�t+/]xݞ��X��Oýp�X��]���Q�~�@,w�f]�D���/U2�	 ��h��y?��Y�XMc�Y��	
'�D0Q{�Hܑ0Zg�W�̂)�c!8:��8;�G{�2fPPA�3&A���D�G5�\�y��a>�@�Q9Y�t��8<��yc�H2��l�衇�u��o)V�:έ,�'�\�Z�g`P>���Mx���� �-���+z��|C�y��}���p��=:�쮽�f��I�1�apI#�uv� 7oC]�,[ȡx�/�������[�:�Ù�p��7�>D��x>�}Z�RWM�`�R�D5
��W@9�G��
�\��"R.���$���	��	a4��嵻5�CdR���U݇_��/��"s.te� ��R� g!ʞ��Úr�%�#�n�:>�mu����%����m�S��Bt�^02`���-��Ƞ� vgz_�@��Ec]��t���14�y��*e��`���F؂#^��='�\j��TNua6���(-{!�#d1)����N�)�K):���5<z�[��y�b����ç߈)o=}��=��tM�g�����&�����(��i ��w?x_�yJۛd�e�9�g���� �x��f�ޕ�_�B�ܽ�p"�d�)���d�w4�G�_��
�H�N�������X���~/%e�xi�h]zi����������{������Q�G�&�����pϡ�p$�~���&�&l��v�Z���[���jg�c���)��$����%���CQ***H���\MPW[xmsH��uS�1t@N�<@��˚)����Z(�3m~)O����tńm�J�� )�c�ѡ3�d����!K��Jo�8����{Kx�w$I[�}Ԇ�M�Nz�Ɛ�wu��	���X0DW��|I�]!&Hf��i�:�w��%᨝�D߂�z�zr��m
���ߢ����~jtœ�6��2@)?��M�7�6�aa#rːoWX?�AŲN��Oқ�V��tYZ6fw�����Z�I%�ޠWfZj��O@3L|B�#Sȯ��%B�S2]�dI\�@G����v(���S.Ћ<��㶮3a'������"��U/:�����F}I�RnC�.Y�����NM����v5�}�m'F��+7X-�	|8R:J�����F����&��f�3%��y���Y��E�zo2�`B 	��Ja�*��1P��ЂA�Y�|�<8-B#X�q,�J�%��$����=�Oӟr|����V<d`�XѰ���nt:��0Q��˰A*��~���� 7ɩ#��ҖL�p�s�����[W�����[��Y�����{E$�,S�#�ؘ�9W�6M�É���^��U���5<KA1�1n�;'�V�����y���]��)v�8�iʟ *���W����y<�t	�B���M�SFO12$�`��_�����W��1��|�o��@�����π�y��RKG���-ZC�;D���P�<�8HUy�x��>*��?�y*�� ��8ǒ���<#�:��eV�*��w\�`
A�[W� �*��-CU�d�g��d���?�h=�T|=l�ld{o;�GϽ>��L�uv��<��WR�/l��,Q��w�� �{��cKC��ݚ9^qe��@����e�R��!.g��L�6��t�O�$b^Fs7�X�X{���TE;x 3����
�-������I�GKrΆ��Cz��F���E�����5��uvVρ ��#� vL �B3i�?S�lU�Rad��D����|�Q<����>�a+� �#��2O���k\���VN�(�qˎA���qd�Ă}��}4�Iy9�e�����.F���1>�S�o�]z'��"�B���M�&�*
bc���3�lr�s��b������� ������}X�ך��U���QEq���BO>����2B���w������G������x�̂^�(�D���gφܞL+}~'��͉�n����JsY���:i� ��9~<"�_3D�w��B��x�s^�~mg�G���7iLU���G\�b�c�E���-`�Y�#������8qXP#�Wj�O-b������|��N�'�is�әo'�L������`�@�0F�6��@�J�|�֊n��J�6�=�,k�?ra�{���]�of�d��6<ү�%h�Al���_��p����}z7�2<���|�##�eA(�JX����K9��q��t�\�?�gh=.�#|��&9���]}{�+���_JM�z���O�Rk��/v���ro��0��̡�}�ܶ�PURo�҆�oG�tef�tX������Jh��)\�xN�p�}yl$�x��m)�Di�mLeHz
t{=�'�M�H+��N�Δw�����.����.�����
�BK�-�$@)֛H"r�, �Wh9ޔ�Z��W��\��l������*���`;�vm�#)Q�j�F�O�Jd٢S%$K����yG����'���	�%��6��V�i���:h��a'���J��6�v�?7�$P��2Zb�;[�`D�;s|G�	2�0��{�������c@W�1�Y��\Ы )�w S��mn��zI��QƩ�g�������%�2,0�(����'ϽE�9Hn�Y�A����;U�����a��-b?�򬄼�0����C�� �b�%A%')4�R[���<�{B�OA�V���:�0���.�};����cJIz�闰�w�JdN9�,f�mi��Y<<E�z��V#e犹�������Ǩ�1L'rL�KE<Np�yUKTs��_`r����ԛ�%�@Q��d$4С��3=%���a���ցəQ,N ᢩ�k�OS���'#�}��d���p���kC�Q,O�s��qR1�E���~�k�w_}#d�c�͟$���w��g!���=K5)�RU�tiu(6?�,į�VU|���v����%�=�Fe�iFL�N��>�1�����k,1��i������?%LƺW�:�}H��2y�������ּ��7R���S��N�܁w��[�E0h~��8j�V�S~�{-�Q����g8�x���bG����9��5�V� ��0F�$]�wo�//�S���ˉ��$Sns33��>K�Xie%�]�aʃ����@��*F��\i�ВTy���a:ή��貂��v��l6]���ܓ �1�_�[�ˌ�]h8��;�W����(�:�纁��|�?M�#�>vo�M��|��y���D8P�c4��?���1�]̗A�"�	ع�l����o�M�k҈T�G�D�J�Y�x�f�!��'9�����$�[��3�f���?�g���@-�y�aV�Շ*�k�L;
H�B��h�t����aז9��~�z���s�⫔qeV�����?�?^�,�GM��[9��r��-����t?�S�����լ��,#K(�i�u�3,}��ޘ��)f��|Y��di����g}��R��Y
x]�sw�*.�L�{���L��8���ca�bR�|��~rAEw��8�ĉ��]g��A(��|ЕH?�+�����{8r,�g�oq�g�H��3�ߧ���u}.<�2�&�.]ǯ<k����D�\�N���
.�7�^�M`C�]���#	2�	��Ofѩ�a��7re�k�À,�%��������x�4�È,S�C��Х����8A�:������n�ƞU���>L)&K����
9�V_��E⫡�ɼ{Ճ�JH�}6�2�A䟥
v-�!I��`�kbރ��ȃ�k��Pl��N��r	i��a�m'�7��i��}�|�W)�-�_�Τl��T�J�ډ�5f�ge<�Ô�$�p��w�0�jxe13�)lQ
>�r��V�- �:+ 4r(�����u>|�T�1q��`�9X�'h�E��6t�X� ����P0�j��y4� ����`��|oTo�8��M�{���FX�O�0�Or>j�=;
�z���}�\����G
��)#��Q���upJ ?�*Nu"� �b�̟����(s�������ƈ�2�~�\�lE�*���Oč"��V�?��@�� C�F���� l`��G�ڈ#���RI��"/O�89���|�JWZM�"'H��6���v=uf���e.�[.AZv����]l�#0��A�!���ĚCNB	bY1n�V�3Bud�ݢ�^$��oLfQ
���oݝL�}�;�$�Ǝ̟�~�8�������E��FE��W(j)��d�d�B���y��jF.f� �8���v	t]�A%}�x'%���.(�a�h�	\�wOܓ�ZGH��F>˅U��
�05��n� ?s�m��pkk32�~��UK{#Z��3����P��L^Z�����O
�z���iK^���BzYX���M8�b���Z���[�a<���X�"�Y��,?m�Wj�:�m8�����`�po���)�T���PErc�s��(�ہT�_�D��
	e�`�0r5M�j.H�u��t����<���oX���t�V�JGe"�|�PjJ�`y�pV���U᩵E u��)���/Ä�pk�4�e�,����k������S�Ȫ�*�|"�Z��ﱛZ�'(�ց����M2�;�>���)ΐ0�v��ZO�C��)�_�`A�1��g���3v3\���Cc�O��A���S����#�[.C��\sN�A�0�WoW��<�~�q� �4F+e�YM*߳k�_�e����cЊ%Ue�B~����r�!9��H%�M=Ȓ��^�#V�� ����.�J�LT/���s�K��1��y�IY����.?�f��h��v�U���|�1j~�6kll�f�K�H��5���qk}u0��>�|SS�ݿ[�&��fw�td�j�q�-�aX8 �_[l���
0�n��}����:����G�!%���-<���R�<(����x��QΒeU�s�~ť����s�����1g���ɮb�Kz�9��&��O` ���޺��ޗgـ{t�3'i9C��sGQN�������~���K⏵��Т{�|���Б_kզN'j�
�Q/ q�I�Z��/�1�wʸ�G���]pe��JBF��� ��Ǒ6Ez��ߪE�7��;�8��&���!�I��൐�7�*Q��g/��r�Å7C�����]���Oj�` �"�����e��$������F�p��7�V�h�����\��9^n���DwϤ09��6f���	�m�.��o,|�]���i�@���E���]�[���^�]�Y`�\\�ȶ�d�T�T������S7�k�Y��[B��D�gjT}q 	c�%h�\a��+�j�b3��X��w�N����[2$�O����-n����}��4��è��P���>��)'M~~у�����z9�����p�����۶I����}a�X������]+|�2����q�[�g�����+\���j�	�7)��l����R��6��f+4Z6g�63h�ŅI$��N2ɎԤ��%�J��ۀ��޹J�5��c��S Y8�3]з��I!�A(�1ݾm�#�S
������(*r�!f}��e�ԇ�\;n�� ENbT�:\tS��k��vE���Wo���`\<B����s�xن����w�c99�z|��i�F~��j�ޠ�#A"�������8{Z�v��FTEYt�,t�,���i�/�q�xYi5<�uO�k$e��_Ip�N��ڥ��.���G]��R�� ���,�M�0�
��-o���jr�HHG��/�@��as�lum�ȫ�ZVMI[���؀��E+W찉N߾[�ͭ�_���#�u�������L���M�������x��O����AWUY�;A�٪3�΀��h$�3>.����Mؽ{#�]�O���(H��
���m6&?��E��H�˿y]�TK	����(,|�AD$|$�$�Y�q��9Q��pv��;����H|Sl��ˍ���ڳ���0�_$�A�@�b���ۑ%�h:As`J"�Ӳch��hw�J�HI�;�T�3���2�JK�fI#DB�#|�y��Z �?�)_����Ϭ@�����m���M�\�r��z�q�f%CM��6�"�E�L$y��b��	��lF�ўE#44�t��Pu�������-\�BG@���Q�C�A�)�	Ĵl4� 6�=�?�����&��������d�d�_n��Q�8x=^-�I�)�*��<�$~��% �Q-���)٭��1��U	5g�=:P��U�T��kՃ*��L����_�
�NT7X�t~ZU,vj�hEM�N�0�LT�}�7*;���6QT]�ûh ��eG��1�K�dVJ��������y���� ")�0�B��^�-������0r�b��MZ��9�b��&��A��@�>���?�m����3l"�h:�CA;i3�<7BI�ٗ��L����. U�&�a$mnVk2�M����ٸC��(�i�ύr����=?t���8���{���W�*��tKė�MBkT�w&���eT�����*�qsQ=��RwT��[!)b?l<��F����6Wʙ�>�q셈�C�)����X�0II�͌� _�������C7DM��|b [���f0���rD������Tpe��gD�ō�T$܀'X`���ȡ!6���7�o�,�q����n�N�B؝���X���B�����d�p���׼��0-���e�\�HG�������9�v����Ve+�#{\B�S�g���t��@d3��(^�G�����|Ϸ�M��[����-&^���|�!��4��G:]F+:�k^e��Gɹ���GE�������%���I`tX�#���#{�&���(W��ލRD+1�5!��o�P0jǾ����͵\<�x���s���:�9,�1Ńdz�r������ �2 �q���3��Ћjn�S�����~���	MvI��Exh����r	mc�iM�~�53��pb�+P/�c-�C�����mW����=AM���G������3k�&#+H=a�yh������b���Wx�\�gf�1>&��E��4%�
每H8i$o�c��j�c�k����@�cs�H��a��޵�K���߇\���μ�r��˯RطQ�ɠ���m�r˱!<ovb��F����Q�<I��o�6���������2⥭7<'�?@�	��0�F��+Nܬ]�M���/"A[b�2<FNx4,t>�8���F�JT� b~˖-��Y9[�~���07�ܹ�sTL�W�)�ߑ b�'0-̨��H(0�����\k
0��E�}P`c���t�~Z�V��[}�̬gꔚ���(�.E��(�����g����ߣ!�X����
;�V˹�^��r\�=��{��]]�3uU6u\u�mKe�E���;b �̉�a�-x���hf����wh���5�g�E4SD���YC��ˡ4r��t#��ɋ��\e�A��=��a��y��L��J}�^�etM���J��T�P__����̔wˡU�'����듬!�錩A������,�����@L�(�{�]A�7[��d=��ka�IB��B��q�eQa�w�B��(�K{G�Q;YLS	�?$�<E)�_Lv����4);�n�gNZ����Y�Ù{M=?�>݌�#����3 f�B����j�	���-�r�.rVߣ����^ч����\� �h_�9����C(Mq���}�NF��q�uC�dV��u�Ŷ��L�励�AC�邋�PD(5pc�A��מwI���x�I�����M��!�V70���H*tY��i��?�-�p�c�r��q�]�����u��I�$뛳?H�ԡ{���S��G�$��u�*v�f������"nd
�S��RÒ����*����K�F�)����d"}�A���*(���z!K֎�0��"��:��?P��h4�� ��k#�̅�7� �<b����\k�{)���Vc�6����Kh�إ�8c����u�>[8ތ{^��/dsw{
����%c��B�5�K�q]��p�,̅ܣ'!w�O�0������m�)��Co�!S�����`���~a���/�'���4�HO0n�?˷�:s4�_�O%��;"_mVVw?�����j,��Q�)��$��M����{�Q��X{,�.6�YK�f
��!f��q�:U���5����ȫ���$`Ξ��V{�����"��w��:��RrE 2�	`>�:D��Um<CaJ�)~����JO�� �K���uoŠ�<l���%��Z�x�f5��=��s(�v��u�N�rA�*{#�)Bx}뿃�O��W[R���f�����8J)���:��y_Rc���)qז��:�/D��?��4?�y����_iؘd#G�F~��$.{�G�k���f���#<�D��K��c>X'ԡ�w%[�\���h�3��Yo�grxm���%7���P�W���e��J�I܏n(�m������������^��$�/�7)jN����������m�}Y�還1�)bh��F^�}T�����Z��L]l�����ȭ���P�S�)��Xkq%���8:r轈s�a�R�S����=�������[= �W�6H�d���W0���Tyl�0��)=s�s�����,��<`o�ـ���9�	v:�`���&im���M�Wx��x�UM.0'.5_Kd/�� ��q��R��f�G�>��δ���:H�.ۍԣT
{���d$��W%�\�F�����_p��i�������t�U�05þW+�qO���}h���&9�'H����"Pj�M���%���7}ntK�����P`���V��~���d�[��4���J�:�������;v�3-�-�����F�g՗��3�jx��qv���)��
c����������z�b����E?�I����t�x�K_@�#����k��=�K!��4�{�Y�[��Ë׈�K�Vy�SOf��5�aE�;8j*j��r��fB�y��x�.�O����h���EU�{��"<�>٣����v��h��l{q��6%��1> gb�rߢ��kc��>E!gg��c�x���n���l�tt��ff��1�L�9t�ir��ᆚ,���,���#��O�;> �,$��~f�ͥ�FjB�*�=�Qj��&P\�|_/w����+uױ=��9�������籺����f�_Q]�u�;����b�X���	�}�^yw�/naڐ�n�qZ�~X����Vg��OW�F\�)�ƃ����8 0�C�9���Iv[$Q%�6b��C�C�s�{�F�9����D��7������ga���v�1Z���C�t�������{�����z��1<�r�]�z���l[e����Ai����\��AO�^�Sg6ǋ!��| �\E�C �+��K"xT__�y,s��H��튽H�Ӣ��;
�ИѨ��9�,��!��@X*�a���Mw�/׮OM���6h\tzH)eRo���>[�J�[6���
�W��:$*-\f�=U�!�H<�k8��5�J^j��iG%�a�����Z��ED�d���	�͕���*�]'ӒtX+�}�H���+���k�K9��5hv�Ԁ��w��(?<P�'�N]L'9g:�g�lV�pv�W�{�_�a�Y<�=Zp�j��P�,���nUzQk_�S]n�a1�5�	�P6�<)�nf����P�C �Nl��Q'��߉�0���^���6R����G���)�y܍��߶��651���c���v3�9RA����IK����.�u4Lˊ����p�	�ٹ2���q�X���Ql�&O���A-Z4v��P��΍���*���Ǌ`��d��w�~+GI2�+?|��Nw$a�D6���!�E����-�k���C|�J�U�������`�<lJ!�J(��́ʡ��]�"$Cq�>��Y�j*�Ӳ�9��I�iUg�&���[� ����R� ���a�)�T�Um�j��DW���楞�b�2y�MC�r�2qg����1ԐbkG�$�b�
bsF���ڻ��T�&Mw�ݹ��4���ӆ8����&a�������x=leS��r!	��л��<{[;{����w\�ɇ�]��p�q����<�h�Wa���a��c�<��̒�Ƥ�#]A�	s�d}]�ϴ/:!j�܂ �NeZI�ņ$'Ǻ"Q@�aG�}pw��z�`/����b��^�^�W��\ׯ��X����tŶ�@^���}S��Rv��q��{�Y�7�f`Δ��!_cק�0[Ru�����E���?n����o-mU��p�I�QD��gm�k�m�h��#�>��y�1H冮0�����TM����m�'�;���.�O��*�x)�z�I��%��ׂ3a���1��Z�6�tJ��$&� V��3�.�7�݇j�b0UQr��
�c8�{������w$&�|aj�|G7x�x$Rщ��m����YP���g:1�E��"�y�w����3�(��֏:w����nF�=���B/���e^�
�����,�#��J��`P��V������+����⬟���n=���GW9����=�V�e�:��<��"���^��M��HV��<��r��/T�ץ7� >]���!�.o8�S���Y)�A�z�C?�S�mM��M�S�c�:"��lפ|.�P�_K��Q&�鍊�%���I�R\����%��F^�F��[4�[�z�kM�)d3V����g��iL��9�,My�rҠ�.xx�%�u�w�����e"E���&���N�Z$��u��Y�'�s+�ǫ����F��g��5��Jm@4��߾���5(&�c�+��һ�0���-ur��r�S���r��*	x�C�Y�e�c�'�d}�RĢ!�>���
��;%���YXa�>W�Z>��c����c��h��z�q ���a	#ū:�S����=8ĥd���hM��F.w<s�[��9ɐ�i,|��)���Ee#hv3�ќ�y)To�B�Q��H�6�`صnZ�Y� 9����l�H<���T/.C;Zԉ�n�V�8�ı������J�ӻ���K&���z�mN�X��j�"j�L�))����~*�#F !�E������JQ\��˗��a��N 9���čJp��y3��T#X~L�*�|�K���_;T����mf��1=���9p�?	 �L�G��^ߵ�0^��/��&,�����a�{|��ħ����ҫ���r��|�p���0v����Ok��*�=y��!MKQ/M�6fL�`�'���٥?@��Uwd�&M!�`_��Ʊ��n�M�~p溜皽 ���uj�W�\��_t⽜����a�P����p����u�ضm��`����O��|����J�bU[��.�yS3��b,<����t�����*�|lK-��t՛�7-����4�h& _`]%f����v���sp������EL��_���	�Q�o����E��X8�L��ۮ�6�)�6W�)�qB�L�9m1*ȅ�m�ǽ(q�
S��d|�j�x����DA3���ʇQ�Y;mk���xN����:B���?2��5������[.���,�D��Nhw��Ӌ�l�����)a8���A��F2v1d�n����3���x�[N;�8k%�6�H�D�[���ՠ�����ǈ�Al ���O����sO�[wX�h~��������Tmw�wT�gRW�\V��rR��W�V��`O苒�U!鬒,�퓁�X}�\��7d�����݈�{&�U��d�ey�Ht�r{Yq�:���cY^��!�I���ŗC�-ؘ�>�i_�iُ�>�� C_.W����=D�oi9�j-�83��3l�6(ڍ�+B橞:�u)zz�mB���:i�5�+`����g����� bɝ��1�E��b�ڻ�
T�a�/�JJ°� EK~�$��H����̜M�����>�g�}t�� ���Ԗ"��+�"R@�2���f��EI��U���Zp�"Mܿ��{X�H�M�aZ�a��iac�m��TQ�����ƹ���@�O�xTɀ7?��_a	�v|�Ʀs��\��-���Z����g����c6t1�)*nJ$��N �T@�H�Fs���i�yԾW3��#�R�X�Bj{��9�WO��Iu�!��0��o���f�k��ܾ���?r~��):�rЃPŐy/���U�Aw֑��.�i��﫚���I)ψ$
3S���(7ཪFhv�5����f�3��k�c����� 2A�JDH�"�WdZ`�$�G^}����K�K�p���(�TՀ->k�J�a>�5U��(M�FGϓq���/���W^k8u��b<�����V�����h�pd:������CS��]8l'�|��� *�ƪSUY�_S��4�]��u�v��"#�>�89#� }H��y^ռC��)ݞ6��������m\p���Y�R�_e�ř/?����笝��GGd��G�U��D���\�/4i5�fø�u�����'!���ԩ��.���������ꡘO�׏b�}�14����;���>�1�ֆQ����)�pt4�!p/�PR���k%o�I�k
)�SC�޲�z�����3v�	z����.�$��zW;�/)(�V��$>�V?5�d	x������g��b��o��W��m?�#c�e����)#�P~N��?����)��4U<s���AZ�d��~_�B��V�A�#n��|����ɶ�=��������d���y7������vJԡL�^�>���FPUq硿&�0�ϼ�(�M�7j!՘4�.��Znp|og/��ѲAB����ѥފcE{�'����Na�}�·G4� ����l���`C>xk��؈�[�ޯa+��ܛah
;5��}]�V|��`$"�?'��W��ԇN&�4�\5f�n���|Z4t��">9�5E!�ƃ�� T�Y��i���=d���PIC���z�ld�;�}MCk�F{�᯿N\`�5��E�>���y���f�Z�[4T_	UؔYg�0:�*:��{6& LT	N�^Eθ�&�A��^�������r'J�?�K�:�rs�*��j�����g�6�5�	��u�{�Z�h'3
G�J�][H�����&���hj������ibfa�ox��<��{�nI(Q�L⻨�eǠ#�I�>H>�<�&_EO��81�N�
[I���tU@��e4��)�W����M����%�p�����u�]b\ˢֻ�g�Tb@#yx��-�&���Р~ �JnF�Q�6T|.�!���r��To��V5���ÿxk0l�1\+h� S��c+`V�,bmE��߲�i���Z=}�yТ-��&�'X�k�X|���vu��q�g.��;J��یJ]�[����iJed���P����Tu
jI�`+��_���A�3�ZX���,+��@dF��F,ny8=�����j�|H�B���2]�C#?�˕����C�C�@�^�b�v<�r��x���_����L�]"���[iy5N��h�q�+�eǅ�Y�|(%�Xe� ��F����gH;�p۴������TL�wYe���C�<�����w��O:k��NU���̫�C��eu��q��-�F�"�����e��N�p��C�V!�Y�u>��O+�wjY5;�\�}`��6h��������-�sAށ�/J�rGIw��4r�٘�,��0��$&�SƍNJ����m�fʒ��eEq �V�4$�ݘ��p�<��ќ�;o���{ՑU�	����Ĳ��z͓X(ڸi��I/��Ade�h0Z%�٪��<	fB��~��1�"}!�TK)D�M��0�1L��}k���&G=�س�c0�(Ż�H�{�CM����&%�Ta�ó��TrW �&��B��qZ��I��Lf?����}���W[�j�l2�4A��7��[�֠1u�����"����f���`���?,���_C�&�^�������IH� ����h��٪	�p�2�'�
��/p ���x��5���j���rz��Uǿ�<����&wmk	�1CD��_����S9ٲ�ʌxcO'�z2�$h���ݢ��A����_j��B���i|�Jb8�-��z�6(x�h�G�
��t.G <aU��0���q$��{t��oj�`��+�8쓛�A���''��r{Μ3��ݸ���z�����a��;�4��[���Y��o]�V��t&�'	F��E�/��z��xcG���(u�2������E���b��F��R�]O�������񑊪o^�c�Z�S��+i��� �z����l�HTi�'ҦEI��Io~;�a���ā�?�;�&��ur���h^?yVt�/��HG�GcYQb	�����U�b��hJ�d��~G��!��<���^R��2�%�E������aﷱ4��/)2/�t`�� �˝�77����{��m��@G���iwg�]y	� ����F���l��k��E�.`0�fT��2�:� �9WG�X-���1�ѷ�l�>�v�N(���@�A�K���������фk�~Ũ�mI@ͼ�M7R(%ۣ�f:��=�r�'��ʥ����'Z({��;���IUkwZ����]���.�.uf�}��k����ngv��j}��OI�w�������������&����,�:h�����B�i�����j,3�rj�;�;u1H9�Q�|���G�

q��Тm��>/�U�r�O��5� ��Řq�ʂR1ޭ$���pg���c19��Ƕ�C���A_�S�#����#�w�P4th**y�-���.���."'RL�#ɶK��K�四"�>Ҥ�z3]��d�Fx��*(B���T��+�(����WJ�ROF��H�b��c#S@9Q��(��u��#��9T�K�|r��j�W���~F@G�`?2��3S'z�a�GJ򭫡�h�J�fZw��6w⥹Sx̔i�;8˚ݟ�"#@�l�� 逳\��y�O@<C�y�DU�n^�)� ��O�W�~���)�8�R�\��_rP�r�ɮ	;-�T֒u��r>�O�ÜEu`�ZE���Y)�ѷ	GݤދN����4t�"�f�@�����` 0��F���5Y	�G�����[�]��zj��"\����!3�l��aL^��r�Š̚�@��9�F��Q���{(�ȇ�D���0�P~�
yZ��e��l�7k����8D�y�S�ǝ!��C���ӆ��E��̼p�^Yd���n���~����cN�] ��1c�Ҁ����s��A`�SK���u��C��g^�|8R?v�WW���v/���I:�bߦ�0|����������v����4c�h�I��s}w,9�_N��x�Ț,��s�H�C�{�U��]җ��SS�Ośpp�;�*��Ӎ��S>�p@P��	�T��h���w�����H��zC�,*3f��,�`M���:�w�F|����] ��S�kg�/�v1XRQ���'�����ҥ�AE�s�H����N��B��h�פ3����S�r�|��] 3�V8�t�K�o�5�0ZRMu�.A&	ʒJ�i��ۣ�v�a�G�-���-`����T�PL����ug�����];֠2�c���7�� (5WuGzu��s�3��1lm��rc�碐
!���y��$a��څ��T���Y ���l\p��t�m(@��E��.m�p,�(��G=���ѻp�^a�������A�|�l�L�r��LGO6���m�ըkI0���.����`� ����]���"d4��W(���Ș�v�M�^�BR��*bK�x ,0�t�f�iBz�F+���{�G�^�<�J�r���i�x5S�C�mޔ�)�`���{-{�Y��.��8}��]�k�f��AiEbK��\����i�fE�YMfV��3ͦ1�������W��z.z���~D�h��fxki��K	����N�zn�#5a��5��<|p=}�|�M#��)SfW����P������&��
��}��=��g�2//AJ���:��h��@���5��:ts�V"��
�Lɏ�M�RA����{�
F��("Q[�PY.�̮ܶ���2.B�K^��%�p��/�K��ܳ��o�o4��cz��A����dtb��N�-/H�����_����������P�2i�{ֱg�us7���{HY�Ce �,ĭG�B�(�8/l}6�_����ab��z��){�os����m9�HW1ޘT=��\��	o��+\?D��y���u��}������ů�w������?u-i��C�q�f?DE7hа_���^$�Y��8��T_ks�d��`����(���h(�	�~����JHE��.AǇl�T�<�0�a)���`���˧��%�	��4A�F�F)��1h�w�Ѵ`��.���k�'��OjO��+�a׀�������.t�������	�M �����o-j�i%J*;���}�b)�54/��-���}4"�q�Q�Z�A�q㚊���ЎHE9�KJ���8DR�0�j�T�x��^�weo�+<�:e��q�E��:;��-be؎DxU�]�ޯ���(S�D�0�]E���e !:�`����.��w�܏!}aI'$�'��ƃ	���z���2"�L����Č�TB�!|�8@�d4�)�I7����I��rbJc҇5���3�iZv���_E���բ�>��r�R��ϜI~�A�e\gj:'�X:b��m�vC �ɡ�)��I�`�d]��]O��R�		˱%������Z,C0�;�<A�@�'��ڗ<�S���obAc���⦐T�?��q^��˶���G� �y�6�s�4 8a@���3B�����z�y%�Q��%֕�=�s�O��yI�s�kP<���z�i����q�j���[�]�<���	g"'�h��$����4~���_��e��Yƶ���!�8�#W�4l��<k�t��r@�.R�0Y
A���,z]֠c3�|����$���؋����BZ���:RB�M�$����/>>�D���OV�I{�!����K��J�ay�B�� ���l:�(T�����r��K\�����?n�O�*�r�dSͩ������c��T�txvz���p�F�:w�!M$�ͽ��x��i�3s����#��=�'Nk��p�M�|�	��q�_=m�#��1���&�g�����y�qG��DB�Ĳ��l�A�/H���$��v����G�����U�CJ���N\4�̓F�kS��<^�o�'�;����M0������ĩ��}��J�������+���Hp���j�:_��[�*z�HÎ�.'�(o�r���T���|*1��&�{����Q~��ǀS��D�OG^�����I��&�"-��#�2Sj���eZ]^к��`t�v��}���owǾ[�2l���$&�TC��z!n\�Ѫ1���qԃ]�,��-Ҕ�kA3>`̜=��<F�����Cszb;E�ZH��^�������-tSooɥ��r��#�O�|�K�b#��d@��~���wMsZvű���Y.VG���UӈUD�RI=�T�P� �І&� ��M��Kx[��Jȯ��ID2�N{x��SW  l��-����cא�>�h����!�C2�ݏ +K�$M�#Wg��	�k-����~���K��-J��8�lh�أ�j(9Z��EةB=W{l�N��j��g���Ǎ��z�!� $�:������7�3d�Հ$ZG9�3���P�hص>$\Q��eWVo&���y����nth���~�	�>"�zRȟ�Pg��N��LR��Ibv:�P%�̨t��bu����r,�Fv#�I��R��-�`�+��{T<���j�95`P��M]2%�e���;i �Y����k�Y�)*ˠ�0�&9M5a�mE �5�����������#�� �}�$�>���XzM�D�� �a d��׿UɚSbc�|b�!�W��WA�2��#��uy6�a��4-2���肭Cg�8�@�����2�aYx�/a��r~9�LzQj.Y�� ^*:hޮ��3�>	iç+Dź�/��5_��Du㻾�nJ�jBN~o�o����P�����Xq�N�����!]%@0��x�,�%6��~f�����4�s1��wt�������{-\����3i/�e6&�º9�K�__�j��+����.��J�g]B�W8���Q2������w�MjMq�p���(�h��	߬%U�T�y�dSm�ci�����K �<n\�0�60γ��sR������F�s��/_q:�\�TV7�~�5���S�\q����t��� Ru�� ��Vq�\��,��I���NQ\])���6Y����}vՋ��;)3\��s��g�`�i�������{���ʍ=�$q���:k���6��f|�#�D6�E����Qu{��H~�ԃo#I��[��vz��}@D3U�M$�8��){����xuG�[]x��'�c����>��H$t�nɴ�x%z����7i{!wdbh�4��6�?w�*�d؍=*��a;o	�F���=���1Z߲i�Y6�عݒy���ю�s�`ܪΆ�_�����P����qd�Zٰ��}�)���炎�����I��ފd���G�VO��(�L4�����8�1\Cv�9X��,�Y�����Ǉ���tN�����jJ��A@��٫!L����81U� ��Kj�)|��3�GԸ%���qC�F,ĊIV�K�#�u���qXɟ�\_����U4����<��JD$Ξ���@x�L�eg1YR��7��Gգ������2�F�i���&f�D�f��H�Xjܦ^��G�#����8E�N����M±~���Y^K>�inЖ��3���3��3�a�ֆf��5Rƺt/��z��kݗ�@qE����D��E:�r���[t�	�G1��c��z.K�]��`�1���d������dK��	OXD��s�0s�j�t���c�L�����A���a2���4Mk�;��K� �J�5��	z���? V�pCU�H�I'�˗{�w��M�|"��f����0��7R�n�'�
�*�4�sɺ���ԂN��E"7�-{1V�%u�Z�@Oy�.wf�D���c�OdN�/+�����ޖ�7>���}���ۀ�"��6�6� ��� ���1�d��i�b�Z\�4��|Uǎb�}�ǖ�iR-��K��Ϧ|���Q�-�Z3���!���j4�ɦ��jj��׸��UiG��;u3����E��U?Z�>��i�#M�wj_D;�=�:��Yf"�u��z$�I�*���V�Gi[��`4�R�|~�ϻ��2��zNw)�C�V>����av�^L�`�텸���B5��i��8:){'�T�����f�������P�ӱw����<M��7HŹ�0���"ypc7�[id����U�� ��4%_�H��e~kcw�|B�� �}��_~[�*3�H�J
<Q��b.q�{��bݛU����9��֞����}�._8el[�A�$����Zs�?4pu�n"�K���xO*����VG�uss�E��{�Y!nT������W�/�e���.
A�cN�g��������gE�/`����;�D��f
j��^�t���<0�UGkFX�᝿9bbr&�㡵J{[�E�����S� �x�H^�`D7�E31O�z�!�Z�@M>���T�W���)���h��a�]n�|&N���lϱ��5�X��￮�J|7*� ��N�9+�옿� ��!a@V�6Xs��{4#@?<!U�o�v�̏6dx��yc��eL@�l�;�?u���:s�Lh$:�;�Ǖ���$�Y<#�.+t'��7�w]�̾&���m�0���0$1hﱬp�Y����;���ꓪ�)[���c�����a�a���>b��|��5�G����ir�e��[���:Pg?:�"]!����l���1�m���l5�,e7�;�":uo�[��o�"f�������	�ܳ4lz�6��Nx͙ho�aea�����`�[Q˸�w^�a��w��� �C�|��[V	�Lڜ�/�x���EZ@��OO�c���R��d��� �A��G(!�����6�+�Vz�ǳ2��P��Hm���?R�H[h':Sҷ��ܶ�K�|
[ɺր#�.��K�^}�����,�jl���^�g��)�~�J�><����k�v���$�����R5�Fe��I됤��~�%���j`wZ��c&�re�:󢔟�eO���I�K�`��g�r�\ñ�o��͆"���k�z!:y�u�n�ok��`�F4)��Yڨ�ʴ歅uMC4�{rV���!�ڳ�{L!2ֽ'�P<!����q�Y�h�fWt��[D.�T|_�0���_��pV-�;�3%T�;��m̀��7��(��n�ɞ��8��}������M-���_��6��u��a��S}�_/�f����o�&5��V|An[O���+�sZq��yc�c��?=���)�c)�[%�)h�4}��+ywq~fӇ��c�������;���ݚRic���U\0n��%�-���q�@�)���Sg�s�����G��՜�9õ@�� t�T7ʂ���n��,.��6g|�ۊ.�Di�D��J_1I|r�?k
D��'&���qU��@v�0&_["q�U�,Հǿ�zFI�F
kMNF�~x� S�����g�,��⚂����ߛH�i����v�A�I�%^l
�5
6��LF�g�0e˯'���^s �v�;᧲:Zבn7X���G��fR	���B�F��qc�Y5�1��G�ֆB�]���!�7��V��ԭ�?�ъ/��%�X�_�o{�V� ��]�?��R݊����3����"Ek,͖�	qq�pK���p��pC�Xa̤��u��fן3�� ����?PO���p\��4��ci#��J�0t;�ҬcZ��{)8T;lT�����D97/�����*U���Ds���^Yd>Ă�%z�r|��b�p�'�zٍD�?�o:�C����v�"P!9�J�u��3|�}1�L�*i����&�<((r�gO���7���dI1	�VC,)ttUT-d! ,�b.�*������2����L�ۡ�<hYVu��*ƃ����jV����|=ͥf	 ���\\ue����s��H�n�K ;��z�D<���$�E� ��.��.�L�A��;y��)#���:�o�&�.U�:���8���%��9�	��ɀT�['���]4~?���l�3�Jv�I��S�&��'S6�[T�q�Țz�����e*�E����5�co�H��]�B$�ر�L�T�b��3{"dB_'�2�������e��^t�9reJG�#s��\�#�R&P��a�6�o�F��!���'b��E_����Z���;�ڳ�1x�tB��+ ԺF�����ΜP��=d���ז� ��͢4��\���\�.P�A�k�b�jԿɌ����^d�=8���c}��,�z}j���F$貃қb�2zՈ �'߿"9�6��Q�Z�1L=�9(��b�^4^͆��)�R9 #o��#'>C��[]n��kVIV)��ӷ�X#��~0�@����/���]M�n@
7��gs 8�=ͨ��
��b���H�_�FPkvX�q�[4�ǥ�]G�Y�8�i�-�<� ���b���u�«l��6kӫc����1Dm܍rf��]��!?0�hT �in��7�:�P�x[:����)ˊ�K3�;-Օ7xF�>^��1�(?9��*�e�ƥ��Iږ�4s)���?ґ\�8�X �A�5?��N��T��(�w��T�����`�يE~��qn��h)"Jg8���&�kO���[����YE�Z�z�#k�Ax'~7S�F�G���A	Xg{�r�>w!��\��	��k��\Ǡ�%�'e���UO�����
OT��@$%��+�o����j� @��[9�o"-�9M�Mp�&�o#��ؐ~V���b� ��t�c'�h�u�'d�R��C��n%h�{_U���R���2FC�u����W�DV��[ä��Z�ٯ"&�(�x�b:�a��+��L"�<�5w af�Oc��av�7���^X3n�C���X�#��zzuo��vs��>B�j	�d�K�'O'�:/� ��~Ag���V�����t젛��0�+�W����)��F�}��g`�*}q�*�L~#�,��>j��Cw�>K`G���QR1���޺3?<~B�����
D�R���4}գ[
����v�lj�}�۔P��\����^� Y"�?w2����cAdq8ds2#�~����J����}�b��IĈȘ0�R�Ⱥ�X[��ro���J�4�KZP|��$LtQ�N�q��L�@;���R�P��FSS��E��r���l��.�W�m�����b��K�r�U�B3R۩w#%7fkf�Ӿ�*oA;�����] I��HS͵�F��w)�����D쓐D�Ia�/�^�pi��.��]I��dm�g)��4&�Xc6j<m^8V7�&��"�%� �(:�UD9����{.���"�����-~�j���Q�Ts�_��b~�0���~J{u|��y�Pn��6��ofF�?:tʢ�#_^�(|7��cW�N�s6XIQ�̧E�g�~�m��\�H�!�U�
� Zv��5���7����F�H�|R���jP渉���w�ue��l��MR>���6�Nla}��D�Ɗ㹋�n�>-�!?�]����P H~}�\b��&@��ɭV?�oA���6n�6PL�Pۑ�4�w�7MY���������Z�7���\r@yN ���rސ��5u/\�3U�m���R3$�r !J��!KZ8ŝ!+�$Ў]	�lDD&������>�c�9�����y��4�����bΕ[��n���Og���IY��C�0�sJ�C��F���䖁s�Xg_Uv��û��}Yƭj�)�DHnVMԴ�k�yG�ﬂґ�7��NQ�����ѮL�y᧱�qҚ�k��-�T@����h��r<♚zZkZ{F��ez�~��� �A���C��|��.mk���Ұ�<�Ż	����JqXB>����#�J78��E��y�:�ۉZ3��@Z7�\��6F@L�l�b��-1C����2�ѺsDC���q�w�Wr}?�j�L��M^�;g�_⃴����ǲ�0 Ǚ"��|��A��.CȔ/��T��J˲m�R�0E��/-��`Of���cpy�إ����nk�^na1�w���&�� *�tzr��R�2m���5���* 
���ʿ�BƿG��)�ͺ�E)�n'�ۭ��V�q��]��K�J9Ax64]���/!�c{�-��>�"I2xZ�wf�E{��]�S�	��2Q��\��=/^h_�#`�J��Ԑ���-��ȟ�^!��'2���; ;�S��qڠ�1Z����cYJ���}�t�غ��]w���9�A߱���~*��aƘZ|�
U5�u$�r�Ȳ�U�����O�}Em�?�nNn��/3�.��ܘ7X�4UeH6� d�4��B.�v.�/��ayv��� r��]��7O�*�/51��+'/0��sI����1�
ɛ�ػ���Df�*	DYc�-�9 Ȧ�z4��j߭����Wճ �����3�aHI8�;�@S��DSlU)�<�c�I���	Z�|��s�.`-��&���t��-*�|a��5�c.JMf�X�(+�KC��#Dc���zv�3�<��}�%�^������s�?x�~�[������\����k���wZy�$�e���l\�H��hS%�zS��1�xG19ym"��q-^��*��Z1�ޒ{#�a�e�D6��#SDTV����~]+B�dz��ʎӭD䂰	�N�I��\�Y����/���Hs�*#�t�CW��Ye��O����#t�!X� ���R�"����UE.�z����5�p�*�H��4��x�`�yuw���'e8N�!÷���2`�!��hP�ݐ��jW��a(��2����%?���J�o�8Ql,E�ʮ�C~&���qc@A�\�Gvo�1���/�J�0{�]R��w�)�a9c�-��܇�u~����M��������J�9�n0��aX�O�[/G5�tKKUWF����e!�uJ�R�4�񇀺���:�|ǿ*6[Θ/�ϸ|�A�w�xۆ,L��@4@��UZ�|�~H�u r���	a绡UUF�����<gos�⨛
~�4vg�7_nˠ������^� �5�x������%A���PܷE]n(~�4��{�����7��"���A
���F�Y��&�C���8ɟ��i���z��IG�'�Z�����*:%����"��cj_7��=�=4ʣ�q�U��&����%c���E�V��A7�Ś�rw=1�R���%�Tp��)�������wCp�����.AZ���q�Kq�4i���_����@�v�h��_hf����q��^�'�k�a�$�����GZ%TR��zr�1�'� fs��u����9�D�!J��у�e��L
)�[ھё�=�DlÞ,Q�����O҆w�6��|�ȱ�X�^:@ȷ�p�b�0�J
4t��ނ���4mUzd?�̖b���Q�@����N�A��8|�t���Vc�&��8��Wz��� ���%ſEnO7�f@�X�	�F	��`%W��
u�;%+�P�KN�*oѝ/�2���O�f@��w����4���?��G�|���8����B�A� י�U�ر1������\��sSzK#�����z}�!q�p0~�b����q��.J�;^<�����&8*�k��u�T-=dZ������}W�.����j[=��zN�)��0�`�y�
���i`�B�&��q�^��u���CpwT~Ä�i;��F)�y��IG����k�4�PA�0�!�gu����r,'ɲ�萰�5%�<�6׍P+�g���'u1I��2���4D-0x�B��#�u�#��1���T�X=��K�����#��b�:3�՛�|s1ܯOz�r�~ާ��s���
��H%���1�;P��M�d�:B�N�c<V�=��ɝ]��j?.�[4���Doܵ�HH/��4�����������8i�<�x�����!�{bkV��lC�ơ�p��tQ� �}��+�2����p��@��K�aK<��V�)��^O�R�
�-89h� \v
���s�A���6��y���[�Ј��& ?!��XssPAQ��aCp���Yx]��?Ma�[���F)k�ǈ���g�=NCN�g��J(¤z�[z�}:����m��G�,dH33u�b@MK
��H1w�(��j�b��N�����j5L���a���묨RX6�i�]X޳P��2�>��tL�,o��_R_h�K*EFZ#�j�|��S't=r��������F"?�2��G�v\y���C˾�r��\���y���.�0�+;G�h��������>��\�Ԣ�#�{k��A�:�9�0�KU[z=���o��'�23ˌ26Z�B��P5f�E �jBi;�#��\ E~�z}�ű��j<-1���М����^��IQ!j��=�뀄��69	�8�: �'~��Y���������}��U�J|?^<���Ajx�?Ø�	Un���?jm��]#�tZ`ÆU<y.�0��Κ��R9̉���e�
��n�[�ɭC�N6�n�?��GU�r	kg����|�^�-pQ���"�{◙�w��/M@G�A���L�{�1����ť����{�{�PƱ�Y�\ Q \$u��y�����NH����3��<�0Iu~c�տ%�1��f��w}�]�9�u7ϧ���O��c��!-�
Z��-}��I��+���i"n�T`�R.=N�tЖ(�Z�4�e!����������F���ubk|i��lx�~ ��]�T��b�Ӌ�H���,<,:���fb5�������q�����gn_����F
��vE�H�rs��{����P�׉�I���V����ã���[�܈��nT�_d�r�r�ںL��o~]�%�����"-�½S�~�d�ԃ�:B-��pM�妒Z"��L��w$#��Q�Tܰ{�k�p�P!rpA���ӂ��	�N<���)	�xg�<����i(� ���A��-��ZDs�ʷ#�Q.X`|� j-��Eu�Z=���j�@=�?k&G���+^(���'�����'���V�I�` 
,�����](�h���B��3>a�~�=4�Us�r��A^�tg�? ����B�Z�̵_W�3�Ƽ�?77��%�H4�����-q�0{mH�b�Z�L]�HhɊt u�jK�O��Ɨvƪ/1p	T�ǿ{��J��Nv@��/ޒ�?�3��̕tn�U~�[q�ע�k�mi|,���=lo�@�f��^WԎ���$-jV=O���ϯœ}����6�����vK5n�3n����k/��?��h{���m����7c�
�$���"Ut�'#ż�b��P#1�44 L0S�'�<[�7#�n�=��X���Y2a��ܒ2���ݢ�peT�iB��B���k$j���=E���f�⮻����M9lU�T�܍��lP� �Ձۖ�o������{9 Կʤ�`�{���T��H<���>�Z���R�ɭg�=Xڙ]�F�"��1�ߍ��'z��Xp鹯�qzW�������8�����$OL?���, ��ݏ��_o�0�8$��C�Gf��0G��R� �ט�6eIr�Η��M�='��:{�X�p���jHb���Z�<tl���
	�`'��a�o!��R��c�;1�-���I-��ס�dO�e�����C�#:0����n&��>>Q!x�^٫�1`?�+h���d��Ъ�W�J��>q<���lTAR�p��.��S�%�e�� \��b�"�K����RZ����{�a� �&s[���Pe��6��Ә���N"�n�>P&�h��b�ҫK���w�	3�_��B	wh/�
�(
}(���諤0����U����7���_t��K_�x$�4ɋ3��>,!��1����H�Ti�񆾵��B��`�f�6�Ob3����xe��t·�}=�io`�F���9����o��b�΅DIH1][*��Z����ͶC�o3a��,��e
7�(�_y�MX��LI�io��^/u���`/�9�Q&7�I��Ma��R䅭t}�a����(v���>���)�H�
�MS�2��4 ��'���HOq�����:_4_>�R�d�V�[��Ed�!�(�^c+k�X�K��?8e�q6vw���u�n����]nv��-��<���W!���=�? T[� ��Ӕ��|7`9����	�����O�jP�+{�+_H��1^�;X�9T�dt���W��MQ�9�߅�*���	r�Ӧ԰
���0]����}��~�u� Χ$L;��|�|$�.R�l�Va��Zu�z���q����V���*r�7rc:Ï0�@�O{����/��!���-�Ak���Dm$1^|���Ԫ֯��#q3�"��O[ؽPB�� ��\h�B�6�;��fsf��<�������� Ă|�L���Y���(���M��ª��?��t���#�ŝ}~�Lҭa�	C�hj,x�E׹\�3�my?߂�2��v�0Q��Ճq5�	]p{7�؟���"�G-�h�U�4['!����QOw���R�+]���qk[w���\:l~��.e0Xe����b�*X�+�_40���`�_�20,./�Y��cb�)Ưŏ'�d}`#͈�F���|�A������mwVU	9�e#��Kk51f����jbD.	Im�ـr�p�4�<2�j�!\�>�EocQdL�0e��."*����;=��t8�x�>�]`������7�D�q�����0�2���c��H�ο�����0���x>1u�U�,Z")]������7�_Ḑ�$IDG�� �<�����ů�Aƶp���\Һ�mp���!��8�7l�R���왨?Ǿ�-��gJ��4��c	L�U���_�	:��V�%���ǰ����:>���朲���gS�w�+��ήM�3Xj~���I���M���Ob6A�ᆳ2:��+���5m��4���Z^?���/Q�#��X�h�"�=���f
�گ���n}X��+��@(G�"V�23�yQ~�*��AeH0�֎��'�S'��.i[4J4�
-Đ��m.sC�y�+�����α
����d
�5yW ���`\�l/̭�Zʮ5X�Q��6�
�k��s�%���yg��5r(��5�!���"��P��b��y��.��Ӛ�X�1)���^��~2!���?�}�����}n�*5��i�uٸ���xE����؏�h���dZ��k�O�54^�&E"v\�z�"�2Hb*d8����Jm�K	�P{�q���^Պ0s��ܐ��e����Gԗ5Y3=�ԩ�$.I%�f;�p��NR��6�P4���JG�^c
5��h*9{I��rQ����Jܠ��5�೼�%�9����?��&�xK�X$_O��>.��/.S���������(��`_o|@rz�
|������Zhj~�V��߽t�����D�N�b��k���9S��<܉;�j��#e�g�w�H�t�x���,��SD7��uLmj��F�J�Zq�ۀ���cV���үTK�U�Q��2�gk���1p�(*z��N-����D�&���< N{��;z���cr*8mS^X�nާ��2eP�.i�z�������ȫq-�"|J � ��}R����=3w��78��?)*K��⣱*�� tJ"z�)5)��1d&�K�</o�)Eg���>85���F��\"��d)�J��*�����s1V4iqI=I%]�L��k��B�f�!����n[�	�����S�cJ�$���@BzU�0N>D�>��yQe�2^c�@�}ϳ�f����+��_2>���!C�#�mg��~��z:�����4A�����]!�z���+�{,�mz�qYC��E�s�U�>����x�;�]�'�K��Tj݁)�x���j�>2=f�A�HT
��F��:�#n�|-�6���m�%� k�q[�YFhm�9)j|,#�n��L�3�,;~{�S���|}�m�Py�^�it�9��D$N|OVKg���Zn�n��g�mWt-B���!�	nLw�ٛ�̷p�,>�p8#��lt�t�k�Z��u1J���l�J�r������F2���[N#2�uO (u�*�g�=��$	A�{�7R<�!�ys�ޓ��dˑ��.P�c��G�m��*�1 y'��J�n>��ƣek�9������+��'�|rt1�j��Chɟ�`jsR�P�,=,�h�`M'�� �E���y��{��ʭ)Z�8z�(��+�/��VI�Gl��Po��
�7	��Gx=k�1u�q�S
n�p��v�Q�q����vćY���H,��dsU}��D��@kY�Ր�����XǍW�h�q���䳕�e<�IڶL�fj�������@J�$L�
-��"j�WXH��o�U���3LQ�|c����v|����Oe�C�/Ȓ�(�~���4`�X_t����`G��2{�[(>����6hc 0O�o��p���/JA��C:G.8T�2Ky��B��_���\h�r�-��//���a��^Ʈ��-��t�#�e�j�����ˍ&N�nP-��"�0;X��L��W���4�Y��z�舷# ��g�Pβ�4@���d628[��'-/i��*;��,L���?[	�McG0����գ̏^��'�M_��S;-�fT�A	K}�-�?���x�l5;��=�������,��BS,�?� &�2*�|H�Ρ�Ր�is�.������&Ċ��8���,��p?��\���Jt�n����K~��#y�x�nB�,K��,{Y!�%��fM�lD6=�ҾL�,�ی'��yI�J�Іl7g8y�3Q�
@�iЭ#{ʈ�/�����|ް�j�]'�<�/�y�`��w�k�Ĩ.��$��u�0��M��+�����BUp�ɢh���%�}�5zb�$�7�n���QŘ�!(7�B&�[�b�1k�>�@�pl�D�A�>��S.<�Oʑj8�}�z�6�T��Xp]��(L�4��X�����GO���b{��bξ�&�9����M�����f��X~�0~Q,:�����{&�+)6<վ��^!2oJ
�|��`��4�u=9c?�L�!Y���K.nv=۵���V/1����,��1f��Ej�#`������(5��,Av,��h��Þ�RsBu z*`���o�L,ؼ|D�P�����!D� i[�?=�W&=x�/�=��'��0���ܹÆS.%��<� #�e��(�t�S��E�4^������Q�C��}^�k�'3>WWLU��[��/��b�Am|����8���cZyo1<
;��<@����+{ǫ)����v�n�[��5�@nч�][m�cK�8����'Vx��i��60�|�)�EΠ��{}�AK�!���)-T&]������e�XK�P� �����gj=˖�����
Q5�-nd& ������i���18DJ���[U���&���vG=�I�X��_���3�\����{+��I�B�I*wˀ�ڃكpV�,s1ZCZ(j�e�6Yy����`1B�)�j#�ED0^��B���5�x�U���c81�|�B�<Q�o�^��&Ц����<nm���KüD��f6}���t= ''%�T"ih�qɯ�Ӌ-82�΅����;�"Ж\\/`y��I�f�M:�ȗ0��f>���Ie��G����m(�m���=�_?���Vu�cL�<��`SrB��a�e���xy�??��Q]ԅn��5���X�[n�h�:7b0n����s��~�H7Uc|���	l���O-J��?/����VZ��U+e�O��*wyY�cc�_�._���kL��3���j�/� k���`�m����+��᜶�o��a�{�3�b�T�������Dr���%�l/�|��E���<�H�Z7`���%�4��m�b�;�[��P�!A*X�y��0qM�BG�˃����m秓�C,��	�i��vv

�0x�{z��:�ۄPZp�����ä߶¾��}3����^jm�lG6�J����Z5sn������.��!��ͯ�ʁvw>��a�����i���N����3`>/y��b���t�}�%�N�dF8��C��C��НԢEx�m^.LeJ^�N%dBF1L�7i����8��s���L�Mq��f��\�T��N�c��E�+F�� ���d��bj�!��-��B&���WLI�K�]�|]������"���_A�۶c	�w������=��V*��4\�nL�nؘҹ�RI�X�.rˮd��D��h�|>Ks�����j���ō�|�=�%e�?�:g�W2l��j�w��0���T�z���ہQ��LD����,k���X�51K)�Iwo�ߧ�/8�q1h��)"l�Q�!����v-n�e�Kn��?)�SWC�\OT�.@���1MS�C-̥BVdW�Nd�:!��9�?�1�#$��,�-��l�UO�E�=���e_P��Z�A:��؋��R��}P��p��W1��\��c�L�5��.�A���M�~����͓�U�4�{q��D%D�y(�J�w�6P��&�a��\�;��)!@X"���?�2S��(��P�������h&����5����)����	B�|wus�m� ����N�82�x~�O�� - �+��\g5�aN�+QN��F�z>��i)a���os;��dI�4l捪ߥp"��߉W:��G�� �o�e�ѕ��e�vo�V�[�����~#�)-�7������̒ ����m��k���PZ�s�slݫ��u���A�|��0����͜�ܬ���ya���1�����A0��,��
���ײ���c*~D����׊m�w�V�'o��*���+�����,�_�w��u�ՀZ����pe��UJ���D�C�{9/�!��v3n�%�)/J�j�Z�	�A�����>7�߷$$�.Wq�?}�:�	J���TE�*& ��Pcq~-�}qx�C��zg'1N����z>������+!�T���d�M>�>e��)�}�V{^���:8`�KFB��������B��R��ҩ)}���o�F����*� ���땢,2*��;�s��N�yR]c����M�Bj�����P���4��垖5<R�lK�@���Y)���]�tC��K����H����9/R�ߓ�H�h��l�`L}�W���̄g�4����2�oDi`�C���q ϘiA"�ޔ8��`��l����6`�m Ch�2@�V�1����B�)�T�Y�EM�(���2X��=x�����<�����#U����a��nhvs��Y����XG��t��M� �5��u޸�Q��؟���̫I4)��j�R���A�t+o�Y�C�:�����t����h$X�1���%�[�<���%��o�����!�`�"�p�i�L?%R���L���K�0x����i��q�ˑ&���D�_'����#�-�h C���ͭ�#�~�Cԟ!>�>JKtt��L�Mf"y��%�'���sZ�ױ�\�t��WV4���1\�����,d�C��#$i�!j����2U�F~���;xu�ʄ^�%&��'��ȞD�Ad_:8���DK+�E��OK`��#�y>|_��.��1\�'X�zd穽	��3>|-��F����w���)z��x�}�6jB�Q�opE�
pk*���Y3�<k�O4s`]�[�.D�@�z���#��!��pUTC�sz���|r��8ZN�%zVǖ�������C>�q;�Va�C.1�_�)�*$�0��z�Xǲ�&�g/�y�^�A�oY)Ε8�O:[D�z3
;Kƍ�Pļ���g��~�.m�����t��_�gw��m�`ՙ�o��q�Bs:���>؝rq�k�S�zX���H�y�xܳ����}���%��B�hS�	�[��y�]l��}_T���o6M@iR��n�@K�rc�n���JR�%na��O�,5�;�!�FK�ju,��<^�'���� r+p^����A�2�B�+�)8��YPs�(י�PIL��l�}�:!zs3Fn��_r?���^I�"%	�K�U༬�PeL��4҅��X@_Mi���Zepښ����T����zr:{Ê������-@�-:�N�t*`��6�T/�Oy[��?ّ�!o;x�:��y�G�;1U��睦'�͂�P����߰�����h~�W�t$i�l+�DDA#�[\F��RQ�)��ڈ�����0��E�Ѝd�=��PC�L����j��A]�j������۱��%�1��c�����X;�*��gV���ҽ��;�wW>*/����h���|E�"%'�y�M�9$/����N��x���)��	��t閠
�D�̰HO5ٻ����_�	�X�����c��(��ou�.�[��)������zP�"lM"̅����ƠN53�u����a��jdVU�K�Cۮ�7��I,#2ܠ]�ah��rd#6��E=�t&���M���E��D�;�v�1P�$��a	����	�!!�s,Aۈ�Վ�̿ c�Hp͛�	�v�oatB���߈u������Z�Z�a�O��4|?y�ی=�� uT�%��>���Wy��9`���Xk!X`!f�����y�����t�A�77v���b&�E�!�ĩ�&x�T�g໖DQ"r6��*y�f���r{���;r:O�*����n�5>�GZw0k��e����<�_Ue�.[[QMF��Am�A�� �w����P	�Oǘ�q��ں��iǚ�4��6=!�!�4��9�Ii��iw����Op�_<E���#��g�9&����I�`��S�i(a�y|��%y�Qa;�������t�<�kk�bî���ýC�J���8�0�������a���]�}Ր])�O����⅜͒���A���=2 r?��� �(}Y$muG��0K�Pޣd��V�ejQhn�8�G<q:P�Lr�j�-B�MM���r�`����M�:U�g�γ#�6�j���O���pɩ��6G��&	�"M�!d��2�7��jB��豼8,��%�K������ ���@�Rzs��T�iZ7{�A5u�iM!�4����I\�0�3�cp���� :b�a��m��j�(�{�ۈ&����e��T�3�fiF�R��&���7�R�ď�U����F�_�J��)���_��)7nۚ�C���>�~4�U��vO�P`�����9���K�Ɖ��2�Y��.�@��4�KJ{ߜ��t��;/�{U+�Q��]�H�Q��AJ�{��B��o�Y,�;�D%'�~�+u�Y�db>��
[^
�+W���
�e�@�#e9_D`���Ρ�VR�~Bܘ��B��̪�2�"�x�Nx���=�P(�����3(��x�N�ŴԺ�q5|���bȩּ"�=efK@��o�F8k���[��.��������:
��f��� ������������?(D5���7󈓴3���I��	������Q�bc���� ��b��;�Y���NJk��-#����[arA�R�GS�:�/!�e�
f�Ƅ��(B�(/�+�q�$���.ۉxZ�}�@�(SLm9�f���u`���P�d����#L|B&��&P`��j����H��5	Mo�����1mR�L��lE���1��+Pь���L��z�w��u��O�K��fv`��I�o-KH&������v��Rpwܲl����OYظ?�@X�� #Gؕ�)�	,��>���(J=�-Ӻ4�cN�e�)9����2|�G��T2�����%�os�����죀8��(uJ��Sw7Wz����6�k�Q��m��
hF�4�ِ 89J=k�O6�!-���'r���a{���9�r��x'�GZ=��]���UB�$�~��"�S�����{ B��Y.�F@D���-M�.a�޿�d�g���vE���Bز�^��	��ꩱh�h��.�D�7�������"��e�y��3���+�'�ue�w�%g��^�&��Y)!�1��~� ���?7U<j��u���A'� ��a�xY�  ��д8�V,뒴� �hMD�(�z~��Y���vq	d�?����O<����&��֚����_���ct�
�ϳ�6|�u��X�z;'@D��h#R�_�]֖@�=���I������Lv`}�����χ�^�k����n���X�����i`�I�+�_/�Q1h��P蟢+��'�阚������)�� �mIRh"E��k4���/���I�s�Z�h^���Ҽ�ֳ�U@�5������-O����a��ss�1��׿� �E����5��M��}Y��pD���~-+B���ǜ�U,�L4F/���#%����6��5���lA���8�v~L���Qy��o�J{��lSq�֪ͥ%=�gX?��Pg<z��3���I�3T�LII�`b��СaP��+�,�B���j���c	�dr��|��Zz���J\~��4� '.��`L�r����c�wY�S�w��4�����i*{���H~z�/�8*����u��Y�����ƺ����5�aF�[�6`qu\g�
�Sor���O�d�Ų����w	Eg�qGξ��G��C7]��� U:�1��)����<��>^�<�K�l�@�h��h)��½o�(�R�6X9ۋ-�Y�H�����5�c/W�X��;W�<e��r/ s*��c��gK���03j��d�H���݅�SF�;�lsg�2�4I�[�G9:'�@���/1�O��<�h}��tXl����x�7�w��S�f+��s�7���B�$5?T��`�;�5��F� e����3�����-���:�Q���W�a:ےBM|�������B��gLAn��Qs�!s�E?��#��bTe�T���m�EZ�dNNC��D�wa,�
U����_d��oQ�����N*5����ի�q��n�4�'zܖ�=����8ʕR0�T�8 �v�*�%9�B!����yQϭ9����T��Fn�w%�>ߴK��O৽��zu����Y����R��2���9�r?�����@��l�p��	'd����)�l��<  Q�B�����B��������iiՙC�<ȉÀ�2��`H���.�M)�Q�yk1��,A�p��,��KzM��ݘ�^����
c��%c��iY�##�c)H�l̍F�^;tZENP��^\d���Vr����ә�Ko���]{�H��ܲ�]�!Y�����^��Thg�Z�r���W�R.��Cw��G���^���h�Z��h��BXa2��7l�ـ{Zň���2"xY��C���*�ѿ)Ok�ZC�w˲x�/0u
�]@�V{GkK�n�K��i�w��F��o�yrbg�e���oRu��V�q����?��S��!U��7Eqs���dv�t<~�,5TI���ږ_q+�A� 8�P5)n7����?5�P�,�BR�.y��i�z��T���ǭpQNC����Y.���c�g1 +q}\9�F��t�	�ҏ�J�Rs�w���,�m���^f������}�K��^2x�&�U�ӵ���ԧ�Շ�����@�����n�/��^��>m�b�9��"�2�k|^4p�*E\ k����Ƅ��a���6`{J�X8�bc[L�jI�dʅq���:�r%�_�d��תӿ�ۖ[L*H��Z��s���iɇ0�S]�DQ2K)uw�/��@
��~��
�eM���*�~�;���M|��z��&�-j����[�\V��T��'�2�Px:��\����'�x*����Gv�	�)q���/�f�S$F�ѹh>��!��/z�e�pr�=_A8�U�
(�g���{A��e��n߆�yA��g��x�:cr+Ч�"�˹�b���/9Kv�`
i�^�m�5t��^Bը�ʷ5q�VQ�>'��$���^��ޑ$�!��ۿ%U�cvB�	�KFЯ<�F��O�F�*�{��n�K�5)s�)��dh^_U�c�7��{�GS�Sp��5�Wb��A ��a?��HY�޾��������,�2R�Z^ϼ˜��Ș���N:��Ǐ-p%j�<���-G�(e�(V��4�㢋l��>@��VtS�y$w#�E��[uJ�m`�.�? �����nrw~ ��)�����'��k�����'�LgÿK.<�ۦ��D��A|yei%N���&D��6a���>�G��<Y$s�M�B�,UD��"�@Qo��L&vY����H��y]rb�^�eV�r�J_�q��|���x�w��A�0d�t1����C�U~E����'â�w�z����
DD����vNҁ���SD�����5)֞"�K"�T�T7j�����zwذ��Ah62Q6�~�@�����m����:����@�S!�؏�<3SDP��zh�F/�,Z<�B�>7)��g��OJC�����xb$a�T����~�s�N���u�f�4��	.��ic?1+�{�EF_~'���$$�d����\�������`������I:�4��;�=a�<�� ��K�w�����H� n��Emn2#�DB�H%% vIĵ���\rh�H�/Ϸ�����Q9U&��*�A'6@K��>)����
�LF^z���ݍ&C�;e
�A��5C=ݗ�j�Ս�wФ�E�dS+?�W+ �3��Fp')Ehv>Xh�!��Uc�͛�za�����i���� �\�99� ��1�U���&Q�5�9ռ�UD�96`^�t�)�]��V�_�q�)���� R����u��WM�I��J�غ?��_t�nò(�} ~'��(�3F3���b{��b��G�U��wW�pњͼr���Y��m<�?r};�Q{#]-�O,���'��.{ .]��}�'<μ�w)��w{CV�
� �,: �"�A�a�uf]�L�8N6�gR��Et�9��E�/��:���A)p/�	�ln����مv��[et)�m�iI��b��k��$�ظ���O�*ZA�H�Y��S�Ȫ��	��	�j�\��O�.�<���z��V��nn�J�©��qa#��w�����<%�����ą�ڇ
���6������fQ�]��?��E ��0AB�e
z�a\�!�o����&9rE4�_�ݢ�^0�3�2`�45�2/��Yͱ�K�n�6v�N1���UF�d�ڷ�K��#���F'�@}�|��=q(>(�D��� ��)l!*�[,��I��rh��#��z��������NS� �;nn�6�1�;,��6A��(1��Ā��F�<�@��f+�~��C\��y�K�U����)r���ߕ8��E��'��oJ���;�yMN�H�36a)�8��֒`�qZ7`�Ts���{�k��	��:b�K�t(���I�,�S"ZE���H�y1�(J��ѝL�iC���*(�����;�8�譣�(����,��9��	M�����DO�)���(�4މ3s�W�x�x���E9����>�@�Y$�^�EkQ�{g<o�8NQ��Q>�-4ag��t��3jC��"h�<��{�r�Fh97^b末2�}�}ki��f�cX�H*�>Oq��*��[_��P��l�"�I�坿s� T&D٦HǗs��z`�(�����E�!͟4&0����A#gק{�bg{���Q���m�F�*�����E^�}��M+F\>���JF_�/ǩ�����U�Ӎ/��Z�L!���/H͔ج�)u���:;���G&���C� &CQ���:�$#x��o���㈾�b��6�ɜ�(�2G~[X������tMm�� i6��\��������4 ��k~���ӂ�荜�>�`8*�W����=�T��4�<O�g$m�ݲ��I�ǋ�L��Mޚn$ ��03���@��:ߘl�Pa�e�jJ�&C��ь��.D�E\�L�[��`c����Ĉ�Žv�����Ȃ.HY\1|��=֚Qx�_��YE�Ip����W$�]Q��� �ZCAZ\`�J��J{ޭw������'�rG�]%��7P�3��)�iQ���{�ѯ�e7+*���&�N\u.����"U J�&�v�B�1.ؚa!��a����C ����fo$O��e��kqJ9�Kc��&w�$j�58zͦPJd<�o �Ђ��۞��1�"?��A6|����R���P�F>�|-�/&��w�)��*8�����H�T՚�8L��>V�,��i�J�C��#�!~�R!����;j���#Cb÷�7�W��=�ҭ�����1��Pw���q)ǒ�O��!��/�yĀ�>`\Q�m��@o��%�2��+��+�T/����'��RK��m���}K���E|�>�ϖa�m���yO�����S+{� 0fZ��EԷ�k[@���'�|8��B9���h���%�K?���3�~_�g��__��x��2�k�Ro�a�(8���b�����?t/~��
mi������'���9��ں�Ea;�n�G)�=�� �v�i�?^���^�WC��٠�T1[\A+D)qPI�����M��\��5).�*.CʥNHܷjBB��b��)��W�.Oul-�gz
}:�!6���� �8�~9���@���_���C�i��1�<��&����㽄�b q�L%iG�
hoK�� 4�[6��3�$[R��u��J�`.�H����fa��7���eFu��?�*�DNz���I�p�w�����D��M?{�8�&љ~j.�y1h/��N$���N������ ������>Ě���xA7��s�3&M�hl�̿4*]�������C��ە,�Jش��6�d���v��f�|�g���N`1�$�'���[*=�1����w�YĶIG(́i�`�FGr��LXR���.[/U;_��=݂س�)#�$jېJ��,�2m��u✞��L�F���4�4��m����?����g�{�J�<�}�n��'�A q�'���ܶ]�|�	���^6��� �M�8�KoX"櫅n���#?�{t}_���l�u���)j,��")f5�H��u�E�{�5&��^�����̖��X�ܕ�b8�RQ|��h���p^��i���-��%8ڻ�?����f6N�9n����S�Go�XW�������('���Ns*m�K�a���Oa��N��G�"���J��t�L��t2�@wI���I��k̞�;�#�d���`{���%�%��ŗz��_��9y3�^�jt>$g����Mč	 �$E��YF���&�B_�k�rta_6R��4b��#��I�s!��n��vp7aE�`x��2�q?J'Z�i1�C��֏�dhʱ~�A̵�퀫��iV��^����̪�]�+)B5%�^�ǜ�$��u(�;�l
�'ͮ�51﬍K�I����G�����#�LK��"�+�˘��vv�߄a�[�[�W_!�5�{�0��f ��ʹ%���Ԗ�l�S��  ���k&����K��p��u^���9i��G����*���oZ����HL�#��r�l.���g�y�G|z�eU{[��TH���i&e,nk���#8���B��48a�Y��'[wL�W�[=L}��F���5�۱�.��)ك�x+�1���Q��J
�DO�-m��� _M�(ZT�93.N�j�I+�d2���;�ܼ��� qҝ�L3D�x��a�L��c�4yHO��ʠ^�ef�6,!t��z��v��� ;����ȯ��~����b��L�	lF#Vr�-	��σ����I�(����z�)��T_���� Ou�y���'��h�c�Ҷ�����=��V;
1Z�t�-eJ�0��:�Y�|�����$��W�������g�P��Q"K�e�e�_.�y��[�t�^ _ƞ�w���`��k*�o�+�?9����t�n�EfS�7?u�Խ*�-�R�wҰHŏ��}E�8�3�#%?&�|�eE��L�#���&���a�wf�T^���DEU�E������a X�Nm�fO�!�J��+P����S�I��*�� �7���uH�VS��+������}���R���)곜Ph���$��w�Rn��q%���d���9S˫T��i^8�k��6_�g��Cmz�W��~�Xѵ'J e|(p"fߊ����-4�g�,�S�������+Q�cZ��;��B9ް_��n�����W��hp�w�SN��zב�j(U���F
9��8�W��S���W��ۋ�Lu^�;�Ȁՙ�s$�Ӡz,J��}@���ݞ�Ez��tE�k�C~~I��w�Hz!Q�m��#��m�`
(��rwc�Np22�5.�#�Q���e!��=KjOmg��=���~^,���ml�w����{Kk��e���pD���.���y$n�Hs�д��۸#j��C7"��{�Sn]q�p-&��Bg�k%�į7z?����X2o]U��3؁���!��c��*�g����K�揉Nr��*���9MR%�#�K�2��}��P��{�m��Ѡ�='�<$�2����Dj�0���\���d�0�N'�������MX�>��afw�=0u��}{�`>s��kP?�(�h���O���)��/1�Ma��.���f�,�.$ ��5b^�3�9�M2|{��R�R�=���Q6���-(�N���2Ud�����M_w�G��j��ei 8N����M,�hD����w�w�g�H�u�m�R$�9|�����4���(ޜ&>�u�ȁ�� 5�R�,G	�ӧ%�H��:H������/4J��I�]M;�}c㫃2�w &e=*�֥�X������~�+��K�Aa����Q�Z�f:�/�w�PYw!Η�a���2 ��i9�M9���;�L���O)T��ʚq��
���./poH��j�n��e?$�&Y�i`�.\I#���Y섽�Sq�-���x}FqsO�C���0!�M�g��Uz�(x�c+�F�3���I���]�? ������>x�xvCS�
9�/*Ҳ�TC�ІX�2IQ�,�[�	�'fu^%�DRlȿ�.�PN��'����ٷ��6��V�سJ	x�?	_�)1���``��p���;��Lr�ep�?͈���jh�:�B&�v�D�o��ܵ�֬}!�u�f�#���VËs��F^$����MY��]���t�B| o��\��l���� ܁+8H���L`�����uH_S���$���kճU�����W��V�W��K4������#�4��B�шW^2�?�-�Y�1F�I��K�I��9�u�L�@�A��RA�;�au-�.|?�e96���jdg�t9g߹k�V;\A607��x��u��]^�pP����sK6(T:FG�gU��O���K�,���(�*T�XRf�@��P�D~��-{r�G�V�lV�U��!l%=NI�s]�!�3�w����������_�Q���~�E���O��x9����s��w�cܦ�+Q�o��܉]��v�*kVU��8n��a&-���'Il���dE4������d�Wc�#g;w_:Y��}��3z[{������y"���M*����8�Y���c��
9T��e�x��H�:Z�?f��^)�_�Z?����\d����a�5`=��]/�v�AR7��Rs���pC�y�7��,���U^�I�� �/i�����!���b&H����1�Y��^�a����~#��8T@�}����ȃ���	:hGv��w�:Z|�BSB�5߯ڦ���}h|%��J�X��(������遇np�_��Ū��4!/�$b�I���R�ڋ�rr�PR� �6�AZc�U�(��ie�~�~�h�X'�-VSO��N�;t1����B��j��+��#�!���n�ԫ��U78���^�7��᭎��{�⠬�e�_�=�9���t��K ������������/b$�#k���>�csf�9Z�s[�|?� �h���q�a@)�-%S���U���O4+������[P��!)��;B�5q���
9\�d���w��TD�hD�pY�U[|R��!���G5T`V�ʙ���$�p�mE7�����[ 	ODK!P���]�T^-&5^l�م���`ϫ��9Ŭ$�b2�N��Ɏq�JXsY�^���^N�u,�������c8����k���ǿ�L��C�1����/��eA���c�[�Za�gH��k�2C��"&�f��K̽��~=�Iv�4���6Ԫ�n�����ij�㠎�E!����4�~��t��b�{� ����J��,`�&@$�:l��rY�L|haw'~��b����k��� ��BE%;����S�}�DS�}���n+(�3�T9��V�~�?����t��霸j�	�"�u�U�D�FmgŚ�K��ª�[E3��l�����f�$I��Y:�Zإǹ�B�<������� �X�EҚ�hv ���EH��Xq��\�J?���ďY�C۪A8�3�8����0�E�8#��cEL�/5���kG�1F�r|i����[��y�< [�Fj�V�1�������~�<��OK2������t�dtj]	o�C�t���lWUR3w?��Ҥ5B��y�-�"l;�O[��rn�Y�Cj�ߢC�H��0��(}j��]ic��/���Rc�f��|-���ẊoJ�Io��Q�PȒ'�$��Z[t�U���5Ph�%��M��e��y��ݝG�;��̜q���Ȑ"�#so_hb�|�5���\�k�W����X��NK�Z����fX����-��Vҵ�.Z�XG�3�d����[4��n�HT�︀t��s�V	�1񿔿��Y4���墠��h|������!Q_�<ĺT�8��"�d�Z�kά$k� �>�Z���g%�������LU8_b���;�=w<X[�jv����^t�ٮ��F����%#����_�z��ql�|QGŚ���Q�Z6��;�w�v���C�Y�0gy]g�Z�}6��$�z������bw�h'��E�؀�4�K��w�*��q�7�H�ƳdbE�䖫C�Y�:�ai�&�����g/���H=��v����|��Ti��ßߘ���a
#�2؟�ZqШ5���'�H4�?�;APLq3s�029��� S�.��� H<.LYӪ�$B!��9"�����<G�A��Z���j����q�ϗ�K&P����|hi�}�^=�� :Hηv=��4��1'��89~L�@�lIݱ�
1gK@j{����Ўw��E,���T��
o������n��ށ���ˌ�ñ��;��9:0�uj�=����GUy�*:
��O<OEzl�y8:��F��p[����������k�s%KvA�X��Ng/��T�'�
�|�H����g^�;j&�(�ȉ��.��r�Ɠ�<&�3cfd�+�q�q�`�_��?8��{�@�T	��ê��ت�G���I�^3�0�1�"ћd�sV<=T�Nq�LֲDm���oGJu�V9���=�����pf��5&'J���6�n��ܘ�`��r���9U:�?c!F�J��V�]檉RHW Í�{�\��Z��΢S\T�TJg���[�~ٞ��@����b 8Bj#D5%�]�6�E��o�8�����ZA��Lj߈���02�	�4#��pŝ>׀jo��)�_z��&׹���<9u+/�5)�s>�ͬD�3�~|�9�g��ڤ��z�)9�?Kh��M�QaK|ǲ�sV>���J�/�a����a�ѝ>2ś,�u�u���Ƽ�� X8Cg�8�gTU���!1����^�w�h�s��f�g�VC�M��q��>�w!~���g%�A�h��*�\%�(�3��pB+�2Z�2��z1�@��$4�x=���dX2[�Tu�4n�^!zԗ�(�~�9c��ߋ
܈��:z������ �9c�`?�ڳ���ʱ���������p��|�J5c�z�1]#�#Ɖ�P�4�z��4��t忐�9gySi��$D{iRXs$�2m�c�7��ۻ��N8c��u�/'��3��a�ֵ�[�H�z�8�?��^�xu9��ऽx%Ԓ��)���`ǭc�A�@��E%�ф�n�C'��E������~���n��)����E�P�W�T��TY�GV�\_�u,�~�}�+�����/����Ev��R%�X�P ���צ/S�ѕ�Q[YMU&�͂P����#!���Y1e����9�*����(�w�F��yI���ʅ��װ��ȁ�*$�P��X��z1��
��-�ȓm�]�7���|�:��_�n�����-��>��Z?�LЎ�;�G%���bz��I�;��	`R���#��T.x��b�֒�]b.s�$.�NJ�dy�jo�l���*��%w"�!�v��j�{=��m(]1����-�0&�@F�K8�x����c3;�2,�"�فe�����:J��Z�=���F�7|��]���+{���]�Jy�P���QI�Zw&�{|y���X�P�S�"�ex[��F΋4�g����k�4{��T�t���yj�xBJ����<������mc�;�ʃ��Ff�q����)��=���U1�Ӱ�}�þ8�-�(:+�egX҆����1���T��\i�<P,&TFi6�ԓ��b��b�� V�Y��|�\�^��H�k���6&�\��P>�pN�G�Ǖhm��f%�E��i���i	n�V��8��nh��Mc�R�.�Y�]]����O��Z���v��5~�1A�y��'ˀ�%}fz_X� �7�p%}����/_��<����t7��G� ��6+�zE����?/���Q��,GE����|З+"�-D&�-d�0.�u���9�}����w������q�����RW�d)ў�u�W���4M*��@i�8��Aìv.no2Fi:��V8"��Ds>����H{��v#(ͻ£�Q9��?W�ߺ����V�-zz�h�Q)�̪�o X]'L���S���}k�}� ;����{��I�)�3?�DN�}��%�����w��B���T��H�N�s�*P��C?
�s��^+@o�d��O�0�[�p6�h맅�2��}/�&����r��bR��Oh]��/�!�{��j���0�.'��`l����Cڬ>�&�T��CG����<Mt�R)6� � ���[tyB'�P��4�}����Q�(��W�&��G�C�+CT�"�b�6E�N�59������'�$p	\E�ԁ��	-�<�� ���_%�@Y�u[[�Z���2��0���;Q�jg�}��A���r���/�<��'�B^I�׊+���P
���E3��b�.�w	����OA�������Z��Y�^27J�X��B�z�AH�yg\�hZ�f�|R�`o{��t ���r4P���yByd	��>���(b��/�.�ij��N!���3m*��7��d��тV����쮇�������`�g�.7�G=�mM8O(9���������Y����������Łb�Nu�pb�L��,����Ƈ`�ڏ�jM���<1pSܕuT#r2���V�`�_�C!M�biiF� �; �A�'����S`�T����8T[x[}��P�u�b��^zi��]��c�h�r���<Rmm�R�Ej��QϿȿ�ut�h=���ͧ�����_²o�#��"{����L�����6ߥ �3��4���_�E]�Tdtj�U�ݦ�⽭Hɺ�++�v�WSD1#�ϱ�,f�՜{j,�����윁��9N�!�f�ҨTHnSF5�0�R:w�T��^��?��n?avs��E���Ҋ�Z�����1��ڷ�JuF��!�`5�y�n���>��q�>r����Q�B���^' =��V\�o\3lg��O���vs,���Ҭ�:�%D�d@�s)�<�8HFSzp�3�N�\/mS��Jf��,�T��,����Et��������{��W� �E��b���N<AhqLA�#.3_4?�f�6'�J>w�(����O�􌝇	��d�q��+�N-��>�����ҫ�͉��󤄺׸��pm�s�K��1>����z�������.-�n?Z噵B+��v�w����K�ñ�p�>}2.M�D&��Y���`OR���G�#���$�Y���2Dm�����˦��~qC�D�]�	E�1��ϭ�?n���G�����f�o��TRf�z�a��.�
�Q 4�����QE)L3��*��85��`k�D��wU��1�oLC%�`4���W~�O��Ҿ4>K϶쑙ؚ�ȵ�_�%��;9��fgp������0�ɴ����%�{�%����mE[�_xY.P�P4�=����̬�rp�&�FܐƋ�U���#�U=v�z����eửr;�����q�)�r�z���a�4m��KL1E��J
AjV�H�ܟ���siA�7��rO-�	�����%�8H8O8���
�Q��9�"�'� ����&Dg�-ָ`�ԋW���I��A�W��pl�$^w0M�i�ke���B$E�ؗWY/
؎ʟ�̾�q:谮s�Bjw��}�:.yB�'P	�}8�����Q�J���{s����2�ȕ�ye��v��}\x�_�x�Y�y�~����$�3�����#�w�df�0܆s.˞b9(���F���˺b`(�u���6����s���{W�j�h��K4+�}'rgB^ǲ���]a�j3�ڨ-�z
�; -�K�A����C.���Oӗ�gC����x��|%:�A�����NDs�k>_�rM�{4m��~Yp��h{�m�(���П ��Y�|:O\�s9R�I0b&��ɍ�,�C���4`4Ih�x�]�'�Mw��S$E�:q��+�X�~Wӂ?b�>a�E�\j�V�����릍�E�:t���#łڍg8� <킥g:܇ˍsf�b�)O�6#�:K��w
��~�@�Zһ�g�Ӓ(Xʎ�Om;����0"{�]��R9�����F��P��*�u��z?���J晌��)Ns�U_�e (���ԣfU�cPN�)a{�X�E��6@��"�*��Ww�Z��>D\O]�[nrs%�&��]��'��O>ڏ�Xvt5B�I�2AO'9+�
���a�S�#&��Q;KOt�8([`	#
-#�v����������Y��:)��s�
�3ZF�=�qs�o���_�^0��E�[1,�������w�G���3���$��hXwVw�ܛ#�#��h۶,�� �aJZ,��2/qOY86���8b�����\0�j6.���`Kb���V�U��G8�!�k�n�E�sD<.-'oF?���Z��.��f��]m��>p�ʪ] 2��=�֎��Ѕc�Ѿ�G�x�'�C�%b���q�ݐ��yd��Z���H���T�ѽ�G�1i�x����n��e�s�n�B���e�lV�����)&z�mp�+/���Pۃ%>���LĿv���u�oO����#�j�Yb�)	��>�<�l��W�������J�g�z������y���v�v���}o�d�7�Eo��	��s�9��1�U@�zu.^�ߛc0����g��L�� �S����6�G���-���+��sĔ@��%�՘����q��%eE���?p�	_&�%�ʵ���/'�#����E�#�A���cH
̹�9�_�/5P��#wM���ƍ���5�M�B�נG(N(���I�k\&��9�F���+U�'�A��n!�4�����zre'U��c����.��)Y�*�$�*[D7/��E0���Z��1���^��6�� ^��I�~6��6E�}�a^��%f�UK�ٰ��
x#x����o��O`����Ay���S��^�U���� �����\̰�Y(U��lJ�!��`L=�_��n+?�-��Y�
���������o4�dZ����0:�RcG�nN���P�#O%���*�F��Wf;��w���}��_R}���Z�!)���\�*�0|�hpq��^���X9v�CSǻ��v������C;�J�ؚ�+�?���}�(�pjP��1@�U��q�]{9�b��N�܀*ρ�n&��8A�t=tX��р���ji�nm�Y���1#�-�����.?����[C��F�d<��Y����2E렉Y@᫳`	9x�2ֻ�g}�}�F����hqjk`���K̥QC�dX
pK��A��>��Qw�**!4Sv�%�3��*��)}n1j�@��?�C��[��c �1�NK���xz75�oK��s_ԏ`���������O�6M,UL�0�D`������䗁��1��X4�"œr�y�q�����$�^�M�E�;F �@7�wVMy�0�p���Y�� =8P�����A��r�!S"�ګ9��o�l��,=�@���+vt����+Z���95�&G�M�)2�.Iv"ɒ�@3�e��r���Q�`�R�i�{H����n��0�@�W};bV�#��ػ2Z6B�0�
�x��Nb��+t��Dxq�I�r�g�b�z$�PaLN2�_������#�Y2{5��So��T���p��<���t'�{����4e���߿*����Ъp����(� >
&i1Ѷ�03&��Y?��5�.���{���g٥�*0�Pz�}&tMF�S��P�m��kR�����s���{9z^���`�	j'���,������vȧ�I��ݔ��r�¾sm���5�����.ʽC���f�)��w�a�!�T���D�x��i��L��	�+�\߹	��5dҁ���E��B�7���-�Hd: �"J�f��Iz��{,�<�tEp��U*�7*K�.�"�E2$"^JE�:�Fo���L�K��>Ʒ�ix����b��|^͒|�ٞ�����_�ߓС��!!CX
��g $�5��	ݮ �$A���W*��'��Y�6N%o�$M��� ��и�H�=�!Z�]!�*Rφ+lW���E.z���ub�9�y����.�S�Q����/����$\��_��
`m���@Sש�KI����v	K�%����)�#�9:��Hٛ��-�?�̂�Нȫ�u��E�+s��R�!�賈�%�=M�X�T|jd��'h����l �}���O��'�U�o=	��!���|��m�'޴dbk��*�IB"�K�ă�Sy.�>K��hr};�볛��V��y����^��V�l�m@�ƙ͋A �%��PK�6����]�3��8�<�6���1J3�3�õQTR��Q�����_�(k��y��*��VИP�QD�|���c��aѵ�g�{��v���CM#3���k<�ڊUL����&�����R�Ӽ@��ʔ$���M��˥ǆ���'u��@T!{�(�<�_������w��r���f��{[�T��b�����/C��:O^t�ӎ�`zW��l�(���@�)	vi�h�l]�0���`t Z�h�a����&<�K۟�o@�"C.��1^R���f�����А	[��.���/����.OVE�7�H��#G��#���y�V��cY�� aRb����c���m>��j��R������򼥡v��}�8��S$�Ɋ�>L�H���F��0���%�sk��@߀9�gGZҟ�Y����ܡ����G���<�3M/�K�W�C������$D��E����w)�V�̢9/�e������W=��e������9��!h���c��-[?�w����R;�rGv3��U��,
�*�܄ކ�*Y�s�^��Mw_�	�|C�gz�b�Pq	�v�k �����
Z'�"k5/C��:������/q綒����?:z^��:�o�ژ牧�ըQ��;	��M��X?Try
�y������}g ʻ(���We�ʓM	�dD���9p�w������$�%\�F�渕o�}$���V!��F���#ZY�ln䆑�:���h�zc#�3~�@��-�]�$N:�ʶ��Z�+��\���@��%����4�NZ�B)Y�aW�4��p�6�Q�HFs������74�N=���ON�z��3�#r=���RqP�������r�%��6e�oS����$�z.�߬[ͶA��0�]���
�%��0��GR���j"?<δ]&J����Z:@49��T��1�(ZTF���LR���}E��N�ZrL�����kP�/�6OF�}���_mJD�����v\|
���xٟ����2W�z֪�ʢ"|����i�~�bDL�B3ǈ��pc��D�O�xGB���7N�A���DI-L�q.R��.�rv��-�<3��b�Xyb��T)�;R	d5��ދ?M>#��Sd�=�G>k�F����.W�BFM�=�����aX�%�>ϡ��+��3��|�B!���,���/�NA�Q.������������%h:���Re-���J��N�zȖm��u�A���\��.�N��r.3����od���6
�a)s�0ypE�������Q�R6���3��}��a� 0�����@��N񙡞��L��p$1�\�@�7�.����["� �?��`
�:i6Y�2���tE�N�EQ�}�L&3y3p��D�2�mc��| ��`�L��oH{�:�8�3�<��%{$�kstC�k��nȘ����^�Y����u�*Vp�ՌA n2r3CZL�uM�zB�.AE�2��.9������&Ie�{I�Sw�aOy�Z����9�{�7Z�FN�S`�:�&_�!�����+hv< /�A�E�����3�Uʶ�Cbvok�NM������r�u�w�����.�Q�az�6$4�[
��ɋZ����V��Zҧȳ�;ݥ_�Y�h�y��aU	�{9���F{`"l�9�C&�}������N"o_�c���ck��)Dg�K<£;`T���j��$w߫��7y�.����o!w�N�"Ŏ*��L���r7=���B"������>vn�Nb^��i]�`���
8��7x��
s��bfhNn������n	�@�!���B�߃�7��R�ar�#u-�<�pk�*��A�b�������Gp��$����V��=��Ѕ��r~'�:L	j�a�0�u��/w���s.f�0���.���E�6E�X~��v:�޽����P�麴Q��� ���w��w�g�^#���W��Ů��E/A5� {���,�X4��Y��6�K����
Z<��]z�Y'VTq�;�����Khs]!��f�Wf��Ӱstŕ��/&}��*#g�����8Ԇ�:X�Y�[,��H*q�j�Wd���V?0>�#��������*���XMz��l'e�Ԇ����I/��SNC�4+ \�yC!ze%�{�!&�qa2��oj֎�鞆d*:=-��B�8g��`���Uh��6s���Ө�B��p��jbъ��mu#�ߞ��޶-���@K ����$��6�J����; �L�i�kʶ?$H�Z��ع}.]g�H�d=��4\/��^�H�DVU��L9�k!�e���\�&ø��FD`P�2��:���9���$���{���]��I�Αq
rX���;}�<�G��Q<h�W\)��MU�K��3����#�4C}� >� H[��� 2�<u�
�I�k:�M�l	ɉ�,g�sI�����;,�;Nkj�5�P\zKK'�΢���c4m3��z�*�]�w�T=��4pG"4�O�����M�&DUN���\�>�$[�-��������<�@�[	�8v`;v؏�]�r��$�s0�5-Y�,;Uc$Ռ�����ɨ���'7cx�> �|�1�$������~��S.��<.��>*r�d�[��)Ek��_�,��xQ�d�6�kW�Z�-wt�(n��t���(�M��0�ܳq��M�n��q�p��_cU���{mҎu��x��9l��S��h�!PQ�l�Z�`ܜ�����MazBH���@%�I�`�׉���2!�H��옜���P�y��1-L1�Q��:cK�A`w&!�@Xv��a���� ��_���v'xΒ�c��y�D�a��=�����:4��#�3��=��ތ׽�
���J�3#��b%��:W�s��4�7n�I�}6�����&�w"���P�L������x��B9m߂�%�|�c:��@E��S�a�w�{ �>������m=Ėn;>��oE��� ���pB��th��d%�QZ���砑ҵ	�/q\��M��|��Κe����-��_Q;�hg�UQ���#+�w�Zu?�"��i>�}ec\���V���d�'*���HY8K�w������+�v��0�s���MP���j� ��@}�rv���u|:Z����p��)Q��бT1i�Ҟ �3%dpO0+σ?�������kΛ��2���/X��Z��P�ɼ��ay�Vea\asKR�1L��ê��2�7�q�$:$d>g+��p�q���܎���-��r��
{eF�Y܂eDs�H�,�\&�j!���+������ۅ{龎�m:���Т5��QGP�+�24��� �`��$��I��ݛ;�5u�-c�^I���"!����~�^�7�f�}ʠ,��C��]��=��4�2�C��N����o�B���:6��w����ٔv�
��{�>���R�TC������Ь<˛�����/Y�`�2��lF3�. 6Bd� �|�j��.nBl�[��J�/��l0pU�^cK?U �NGW=��;p�_�}�)5V�$p��lY&��v���U'a~�hF&ݯ���YN�����j���d
߽�~��+�nZ� ��7�$X��Z��q���x��G�I��45:$y�i���!ix��@Z�`�6B2���+��AGkB�������UrqY��l���̏�M�(���r���=�J���׻+���sAEH�=R��]�K5����R؇�Z��Vp:����(RV�ӊ��m5��o1�f=��"���~���!�_6n2n����[	-����T:/`��I�d{������+ĸ����w���m ���c�nD���%�-�{+��Sa�X���*iR�w`��]��	c߻0�.6�V����E���.ⵒ1t�!b��K�ί3����?��@�0e���b�A�� �Dx�E��B���-�֯X<7jE��f�إ:�
d$R�h,�KPn�%��`#/Z�j3���Kr�2%(q��m܇�Ĕ��F�
�E���
5pD��Iο'��h��h,F����o)StU!q���tϝe�����19r'Q�H�-�[[CmR�W/CjJ��T�¬�/Nn0��!1A��<8t�ګ��r�p�x��v��[��׭��$�c+,��מ2����7RR�M'�g'H��a�AS�  ���Q�v�I��v�W4�͜�y�5�S�dcg,���KA���fWM�q��*��Ů�y0[��5��B��-�{�9c�'�"A*��ܿ"M�M�Y���.�l�{�j�Z��mZ��[l���s�A��8Q��K��>r��YOfn�:�Zd&B��}`�'���<�������V��S�)X�C�}Uh5X��h���E
��F��l5T\�������C��p��LL�G�`KZ�R굊�\&���I{�>�Lq��9:���M�C@iE���x���S6cd4;�P����������3���ջ�.�<���u{J%�[&��9�U�o���d�'���n�t+��
V�x�L�l�����\�n�.�I`ǉ錁_�����P�m}���8�0�Cj�Z6���Rg��X�uwҶb�k�
&}�AdCbxfy��:
����^��R�w�D2�����$��)���	���D�r���l�oܸъ��y�#�(Qx.z�@bh�7���+����e7K�\���DMuAm/�R�+7}���q���pԷ�tBʧȜ�~d!�]����p�Y4)Ҽ��Ցx�j�q���J`��k���]�&c��h�
�h��j�X�Q=P,��۹˱4ϢA�*�
AU�.�;�f��|}t�Տ�����J~�#yN�E�M 6ʽa(h�o	�)�o�]៦W�l�g���6�uȫ�͟����7�wB�A�O����uXh�d��ߧZ��WD�$���4;ؚĬ�$��f���B`A��zI`հ\o9�w0����w����`���]�
H�)J2�bq��R*2��m��$)�.%�=�%�mI�����NBWX�z:�P�ս�o���FF誺� 
�?Dˣ��ѥ�Ķ�X��b�:/���d�ZB�7���|��#7�P��/(J���*y�����um�7�E
N���l��)��7\�� V~rki=�f�(P�0�qkN�Px�m@mb8(��H���&�:	�I�RB�vc!�L��PgS[�PjI����eW{1�	�G�!�K�u�AQZu�����a���2��r����_��B��G�V���Gi<;�&�&�_(���C�\�#=������`B(�����l����!��w�YC$#m�}�5#5�'��O����3U����M�j� tՄB$��Slŵ�leTݾEC�S�]�����)�b[��ǚv��Y��)h���(,�Ve�@(]P����*߳�c]����`{#4�"$�pmRش���S�����O���6���B�f�����B-�Cd�)���eF3aS�Yp�0�VM2�eM��g%�`�� 9KC�k�܌�T�(/�S�!c� �{�xvu�ۼU���5"�u�P��#��nǖW���rYs#4�=86H�z�5���j�w@�co�x[���Zx�grо�b�hlv�Y�-���G+���-�&$�Q0�J��?B��M��2�Z�]�̇ʴ��8����ȱ�P�oѥN�)�#Sy���I�����Ƞ�	ӚǓZе��%��!����2�5Qe<��2n���tݳ���(/AD���<K�DKnA��O	��N��B�d��J�"}�u���!��%J���#�K�@����<�b�n�(�
��§���D�1��!�%f��B:����)W\�[���kk]%��J�ӦB�)�1f<�	����3VGќ̇�F��=��&�Q�zIAo�C�JG��ӑA;{U�[����7Pc�&3��+���!��j���NA�Qa�:�bx��!I��{یh��x��#�P��?(yQ�=��9���tS���?�/o����_�,�'�~|�5�ֿP�Bh��y�h5��d�(��x끠��p7��m�Kk@�oYȬ��#���"�c�$�1�h ,M�3K'��*����>:O9��$���O8���[�󲅑�����W��d��dG�v�	�X����@���+wl1�Ԍ"{�+�*��|t�4Ft7t��0c�ԝ��U�F�;_���Q��WF!)���p�S��8�����
�4�Fv���0����_�<���M>�IX29�!���W{�op��gm��^�X	#޴���Y�MD݄����l��'L�?���4�CFȗfn�<a���)҉n���:0z�c���O���H��Ӷs�x|��,b��HF p�W�LtZ�2^x ���ǝ��OzE�;f.	�z��qWW�6f�%$A6��[:��c��#��{	R)�׍����]�F!|t�)������rܠ���O�p�tK/��ب"�0��޻��_��g�;�u�q���sI�7�\�wO��+������� ��'���l�<2)�׫�ǵ�1��R�ؕ.Ѭ�����N'�C�V��;�{o�.�6$N�$�mvĬ���qF��Y 6A����a1�)��� ��D���6G�]0}��U]��m�);Bh=��Xt�����3&���הd�}�lnG�㪔!Wюs����vu,�ɒx�S��~i���v��;f̱��=��+�&y�:��*���-ulI@��f�Tr��`��V����4�>����
����ӝ0�L	+iA� Ce�B���z�o	fߣ<�Q�hɷ( O�v�ߖ�)-�!�A�iR(v�����.U@'�͙��4'x�����9��Sצ���3��P���i���̲I�#Б��M�DI|id����3���K��k��]w`�K��֫�z�}�)C���Bc��C7TK��R���!�54&�؏�{�Wd��H/ބM��t>:l	I��bW�(��PC�pd�my>��K��X��48��΋(yo)��sOc����g����Ժ�W�� ���$vJ���')vs���w.�v�&������č�g~8���!��5����Z�obu�ۻ���Sd T�{@4		�9]�|1��j1�KOHO��(?�k��v�n��t��PB���,��0<�$At��D@�����pC| a��G�M6�R?���yS��îLA'�2,�?d�k2�B���o��Ɇ����?��]���iߴ�� ��a����B3���]H�Jk�֌�&�6��o>8F	H��o�E�n�
�Y4:"z"EP_����ӓ��{�IG|t�-SFy!A�D��jg�̀�mo�(�ޠ��F3#��X>+IЛZo�����������$<�X�ƶ�+��;�ǒ=crz��}�zM�Wͧ�s��+b]WH�/n�������l(+ცq��KM��%k��X�\�^a�1�S�}ʊ�.i�-La���k��?eo�E�:�gn�iϫ��@땟 �GeD�>�\,�~�x��D^V�����j��ɯ$O;8ܠ�[�.~�,��/���b��.�{K�O���-r@o������s�$8U�j؟�����%4�z��QS�nP[i�]}�u�?a��-I�B���o�_���1�/r�Zix%WP�=���س����*/���Xs�_#��ߡ�p���^mU���{��o*$�B<��n���V�:|&�I��T�X��1�q��E��Ы�D�U�����g௏���IK*Teo���s��g�e�T�,7s�D?B�-����l��ͯ0���T[�^U��	���UJ ��c9)���9"O:D�'�� GG�P�O&���p�[��9^>��B��=D"C��D��~�<��2b$��gտ7��/��≗�BP���㷾��x޹ Z�?�i��
5�
my�)b;���?2k���'˺��=5�۞��ef��W ��������W`�(^ꂞ�A�@�m}�)�|@9��ຠ�߀���#��)��[K������a��Y�m�p\}�0���`;w�&kbl�4D�(9
i�	���J�_�p�U�u�����Oe���z��*�RGK$�����'���x�H����qZ�60,���*4�I�^*K/L�a`m���s��lE=���a83��º;��)j��
Ϟ����*��������Q��ԢQ���[�f�fhh��ƨ}]��(jV"��,3) *�kS1�&k.m�^�����e�݋��Y�Ψ�B�������ݳ!��d�:@��������p��
H𵷆�{̩�^���o���M�c�j�����/XV��e�`�̊�=����1�+�Q�Q���5�|Y�G�7�wo�E!�Ôg?��P�>c�ծ��q8�pG
{��3Q
g(�@�����*�Yj�Gld��a�(��*w��g�ww�)#AJ8� ���vC`Z�gYE�BbP����W����5����,k1(t۳��XL��n��K��-D��JHq�N��>j3�pq-�^��s�:�"���3$-�tdXi�T�����*GqF��n������?[�����t�8�$�9ɢ>w������T��V
j1�Ȇ�SH�`��P3ɒ�l��^�ʋ�-��	2���b��j�A0�6H>I�h$rrI��CQ�"���=b3I7��W��� �c:�����C�~rA��h��!6������T9v��G8p�#������t[۝�����+�3�+`� VdT7��Dj�&�Ywz�v�݂a��ƗJ3qz�m�C,�cY���f�]1���@s>��+�v��.���4��S����n�`�w��Ǎ[�wT�xX�q��'Vp�y����D�'��S�:.�*C]zݫ/sX����P�x3mK���!���(�����9V�P��F�2�}������6�%%����Pɱ50�K�杼&6�?��P�0�}�St��W�1|,aO"S��r�* �t<�Y�D�#��� �F���d�ۭ)\���Fq:f>���Q4`�ZI+]M�N��@䊙`-O����%3vL�EZ8%�x4w��S�uX�9׼�AKYƑ�Mi�DZ3��/H�ؒյ�߫z�{��D��k��T�G�ڡB[�W�e����|9���� �t�\ c��O�@��/
A�����S;9������X1A���5�TMl�ë��rd���	^����Q����~N ���g{�m���}���2�Z	������R���y��|�k�G����Y��ak�h�,A�ÿ�85��Y��7N���9k��P���l�jt������JT�*�R����?1�ۀ�����Nr����<���g� �=��� �c�0��^�45}zV�ڠ5VY�Qy$���wV�$����"�K�(J��ع>�qj�.^I�����_[%l���q��_~�G�8�1���R�W��VF��.}%�+�	^��O?h��#Iv�L������o6H�V��5�$NR��h�Kf8��d���2u�}㊐=�(ʚ�#T�:i;�.��Έ�[����6�����=����zN6�<fy�ʟ}yV��? SE�Y�_�`JSrBA��U��\R�֑��ؕN�B�"���3�H=l}f�'�� �pU�E�1k�ݓ'��<������ښ�?D�NRw(�&8*/9�/B�g�w���%m���7+�l�� #��%�G�0<"lJ	�*��|<2n��+��;��9{(ci�߈!���8;�D��^��ϗ��*x��xV���yxל\���e�D��&oh���*�#�^��?�n�m�&F���c��ݦ�t����앥���%�E^p��!����WV~K��5e��t�t<�U���<��B�P�Q_?�T[�n̿��ld��������.�kM'���3{��t�]mvv��]lޭ۔f���{ �v���%�bG���_�;�T�rY�X�'���j;]�:��\
�fȝ̖�l�V����̌i�`2���ѻݴ�E�\���j{�6��!L��a�o���a߁~z�܆�y���/������z'����*�	��j3�%�&����ja��a���������А��99��wkRm!�5�b�z1�Y�J����J�ɨ��>���S��i'ד>�sj3��5��o���^����h�=��	26�uNq�|瀦�́�/��|���^��v��-��;��N��u[S�[�;�[�Aqٷ�n6���;~u[��1���(=L�0�bS���|
�/�<�o�!XK�I2�ˉi[�o�p9��'J�o��GD��*��:��Ə$ȵ�3��[����G������S����H�2���)=�����j��-81���R���������ل���$Ԁ��]h�shh��"�n$��Uo`�J�~[�fN-�0��袺?�O=�1��|�����>�W��2{�n���DqWx�T�R�xˑ(���r�4�k^�,�uf�7[+�%�5�L/<�=C��G9K�X�d���P��}8�&����P �"�/$E��ܨ�N'����./|d �V��Vqcp�쮼�����LŖ���'�.;���M�2+�:y�B4^�+N6�3su�(g3�y��1eK�KI�W�ڶ�2�'�ϯ3Ʒi$_V����YD�(Q^��	��`��Nh\�g��9�bףRLU*��H^��D��X3��UF�&��	� 8��h���3Q '���SȚ��<�*�t�� ��{�r�L�[����o���^1�r�[�����Ӆ�_}Lh�}�]��t�A0� և����|5#����c��FV
[�����S\+�M�����CQ�Z��#fɎ���,��:Sk��#����dចl��8'!)$�d��-�p���3�E/\�)��2��Yg�`%�f��0o7ݚQ�!#��v����9�� Ҕ��c]�ꍽ��8X��P
&t���'�=M�n�7ڣ9����ȍ�#J�J)Gsy��X���{��FN?�E4^�+=���R��^�h���y��CD8��a�~���G#70x ��wz�O.��-+�?�gX�Ƕ���l#~��x��|�|�ͩ�"M�m��<��{�1����TJ�g�VB<��?"�@�+����L�}y���	�ު���`�PQ�d�r'�P��w�' p�=�D[[�}]ʨ�t���~t�Eid������G�3k��!Yt�w4�g�Ɖ�W�G'��*�B�8�+v?GB`�Nϐ]�^�Yx��������].ꔲ���M�z��x�%|ۆ�1�┨��� ��ҭ�e��$�]�޵�_!��έз��q�Cv�s�k{��ٖI��MX&���V�U�4y$׏���𷂓�+�H����8�T����}��!��ȴ�#�b��
DL�D�T��^<V�}�W�(�%`R4 GXS�d���&h��`�����]""Y��Z>��?ؾ�]��[��:t٦�����3��֑��Sy0��)�&�y��-'j��s*m�X�NE���37)����[D���hw!�M�9u��	��g<���=��]g�T�����E�p�7q��Ʈ��F�2�����c!_d�U_�q�K���@�Uc\�q���$/R�@��5�t	7a��E�8�t��lCX�sy"ɇ�esV��!�=�w*���sR�6��R����<��Ω6Fܸ~p��y�J_@j�>�����g3rQ|-�;�e`79�7:ǉ������~"'V���5��Xr��� ���<�^Sfǔ�R 0�d�T�룿��b��f�P[�7��g���Q��n/��l��5<�*�Ænu�(C���Vȼ���Xl�P����嵔�7&=�\�oU��֛fi�*�o*�� �')� �YM�e@�MQQȅcSd����I���x��L�ቖ���E;��u){���)Z�6��~|���	���$\+�^AD��ڕ�LFbTאD��x���QXcO�^H ەz^��eB5e��+<D4��7��V]�~�	���}y�;ӎt��T�ooS,>I�/W�����?�>vw_KZi��g.������oǜ�m���Tã�3Onsx,gf�jwyEh�������Nzj�c��_�����.;��@�E���N ��������ц�������|� \�^M�;\�z��lጸ4�5��E�$�-Xv:uwQ�d���ȶ��x�_�@(���6��mo�v�L���7���f��T?Dܕ]����NJ?���pæ�D��:��Y{��Eؚ����]�\+�k	9�gn.�����g.����q���v�md�Y�iX	u� G�}{E�c�P�g��G��� -���{��<M�m���y���l�JP�lt0��06���Bp���;MhZ,�S��X!�Nc���6b�@��s\q<bBo+�>���ׄ����!���ӵT��4WȄ��r�����4�&�{1�h�W�u�\kh[@�f@���-�Q��yv��T��`ϰ�􂖳l(���v!���'̕ݓ�W��3,�Z�2������ݷm�5�( ���yy�!����xR�Đ�W�4���=�Jc�Nn���PE�~2o-8VU��
'�*��½Sn�����
<p-��$���꒣����*/�ή�t�_�.���]�x��7~�ީD�S�J�T����<�ً҅���bh��O{�y��k����A���Jp�+^���9FHޟĦ �z쿽��^�{s�ݾ�����iJ�V�,v�9������r����`"bYrW���"xq� 
��ĳV<�TƬ��x*�]mk!�ʴ��g���[[�ޖ	q�B
���W�Ap�V>sb ;x�t>ҋ+h�ޔ2�t{����z-"��5�&연�VsɷΡ39�0
P��[��v3�{)����]�2���K�ĮҎ�w����}v N&���U�-�+�D��tb�ky�%.7��T��fm���{X�k ���
M�-���U�鰇�:��}h���z��L�IֳcH� �iK�}���\�W�4��Xc1�q�i	=�t����4�%��|`+yb�?�^����Ű��j��~����ځKi�m���©��^����Zx����[\��S1��ܻ��H�F����IS�>��L��6�p�6a_l-Bϟ��"����0쁁p>�4��O�N�`G���C�}0���}2����C뢸����|��7�Y��s�gά��c|(��7&=^񅊐�(A8����D�LX2���)�u|�$v�r�6����:�Ʒn_� ���`��`J�d7�������0��Ř�)�{��ג��Dv�d�$7�\�	�n<���t{R�	%��m�t�C����Ê�T\\��o�C���kṚ��p�����V-�y"a'��YY|E�"m�� ʩL���77:�-׆6<<�g��H�v%���{��J<hm|�5��o#���� |\E �R�S��m��
^�h �!-���Yy73�ֶܗS���Q���N~;�t�Q�$�ќ,�h\M��ķ�s�1s7�l_>K�[�S�{��X/�M���ʹ=s���̊�!{O��zul/��/�mlf	�y����I���W.¢�Cγ!:��}����"�mq�l���'�t7�A��$u�-����sOר���e���k�@�mJ�����}�,�/Ln'UQ�!�/��>���k����۸�4�a��0m�t�,$��^��q�,hd�>�/�������2�ô%�X�V���7*�
�K��M��\���Xl�����!�����
�g�><��|�i�rpǞ7����SzFk~��49�5n�z��8+��W����TrF���i��b�M'�����~Ap~�{��^�6V[�܏CT�K�t*�z|Mb���^r6�|��ʻ���R�'�himYc>;@�� ����Q-�k4�F�A y���q�?�!G���kpk��8�[�/I"�(pd��
kYH�0�`3!w�F��#��
��_i�hF�G��;O/YL״;�d�IZ�fJ����(*N�
P>Q{끻i�w_�F	|+�l���nf�1�����`&+���r�F�D�ES��_��_L��Hi͂m�ru}F�r٬h;�4� w��ߪtqc-��X|�j���<[#	Wdw�}*��-�	rAr9��?=�LU��{��z͹�����qZ�u��ҥG,�UY֊�o�r�/@�Ƨ�.ֱzN�mD��j�U��2V-�~��ە�ީ�,^u����~���t,T�D9V��Ꜫ��e�nm�~�|���?�5N�*A싓	o�B;�v�]�p��m��X�Gc,����� 
/3Ʊ� �Z�hr�ّ�f����)��r�˦�)���L��]�nq`��сm`�2G�7Gta�p���|\������sخd�g}�h��˪���Cd4!ryxI�^̾���}�@�f�M�6�^֭�7���Π�5�s�pDҤ�^믕�|ށg� �
�P�e���x�;����{ےP�5�Jʇ,��,.��(�XH�\�%Z��8��|jL�:P�&E?�]��U������<_�(؍����GAAחD��(�Q*^Ql���v���Ni�Q�K�|{��^eتm��B{rK�x''�k��Q�j�J�H>��#U�a��L(K�9��i��\⁼=s���^@�{P�R0p�_��W���m�c^������L4ӞQN��eu���	aV��&o~q�q��Y%�yL����8��?����-�7� H�N+�#�=g*[�h���Z�,F%^mO��$��\�"?�l��#�O��)�׾����HW�/6sw-�7�2�&�j}7Ў���U>�ewt=��3�mג���a���t��%�ߑA�$O��b0B���f��Y�@��\%��.@~9�T�s\�s'G��ݦ��<|�6s�p{#�>�a�:&y�?�!K��Ez��yw<)G���`;��R�3�O����͸����4�ah��+2R�Y�Rp3B#�M�C�hd� �U�$D�*���bh�J%HoO�J� ž��̈3������^�D��M!�c%�l&!�x`��2���iwN��
�~>H����)K\Pa�{s�϶~�=�1��YV�h-zc���	�s���p�w��rx�ô�~̑R�'-~jt��1���lr#�N��UY�L���U�97����lA~^l̢\���f�@Ea��j4)� �q���0�{Q x�ȝ�w��
P[��hId��]F����-79�������?��+�{��קw8{�?;�pM�ɰ��=w�]���L\�r��]C��%��AC�<c n�#�[VlQ
�
-����@':Qc�#\�򈸹��["��I.��P��]�(EP6��	w
7����s3c���dQ���h5�(��pn!'Q��o�IVJGK��֌��-�%���7T�N����ﵩ���G�o{��4��-��W���#�W#�Y<��kr|���tBU}�\�)�|�@���LUfe�јm+L�yj#�j�aO�5߁�����9Z�����#HTYف[>�W�!i<C���9~��b�iQ��0Etb&��E)�HS�
s(3�׶+⬰65"n1���{ܒ䍲��|�/�̰t�v(@��*��<?x�-�O	��2Wx2�U/�vfd� x|�)��j)
�=H���)�t҂mv�n����4��({w�4Sa��na���V0} v!���# ,�͡<-nC�l����8-1�Δ�x����8�����W�1����޳���
^C�vM�uh�F���M��0��ʊ�Ūe��ѵ�I)��6'ۈ�j-�o�^��;ש*ڑ����3ŉDW��&l�w�&v��$�����WNV�t�LT3��p �$�1�H]�(o`e�u�����<l�c���}�i�(��XV��'��QY���Q*��3*�یM���㓞(�o#ZIդ9����C/~���	;���*8��Ү69��y�JTޒ*>#�"�T�>��Y����
��[�~,�-'6�de�6eu��+I����E!&�;$}�6l�s�6a��X����ZK���jD4y���^b��դ�I�[����� <�-h΋�hA��An-�1��݃�T�I�s�jX�;C�$�n���'�1��v	�7��P	y5��j�Ƞ�e�T�l��&�ɝW�)�J�������zxU	Ԓ���&�Y���r9� �3uI��Jb���֔3UT5��⏫j���;v�P
F:���i���q>���A�4{I�u��p����9���"π���ヽ�S�2�+��z�xf�&��Á'ku�&���:׽�]��n������W�uޫ/�����i�d��m3��6f}(��m��J�}�7+�V���S��eC��E�/�K�]��bB�p��la�M�1�%N�j���[���.m����e�_q����H���p����lb������|j����\�̑(IJ���Dc�2�P��{ ՟���%j����9z����6:��a��ɕ,}��R��x� �srlf�I�Dߗ	c�OZ�_l� ~���X���Y�ډ�o��G�h	�v '1�Y��Ynf��ѥA�0��>ʽ������[�i�#����޵b6*f� �z�jԓ`���w˭��쯌�nlK����YoY��Z�$و���o�rDY	�E��4O11n�/۪��Y�&�����E,��Kn�����4�)�7��[P�2�j/X�ۮq�����ہer�h������K���֛x�Jx�*�z(@B�/���C��lM�ǜ!��8����ʡ�BM�K`��g���Sb�_�^�����aB�e���3�����M:<�|��)<�%^J�.�P��T7��2π�H#r$l���������Yd�����'�~�>�1����*+�k8�*t�	���Cd8DIN���MǤ�TWg���\v�0�d8JA��x�%#)��M�tڊF��fՍ��AI
��ֳ��N�������	ۘ`�����.�#�j	'9��0E��"���s��`�c�xM�U&(��y�������|���	��T�wyU�v���7B;��.�PFq�0�:�H�wA!��ƙ��(��ш���d�����m��UwvhT�P�@h��^\ �����*���<Rj�lPiB��7xNzB�`Ɏ�.���iU��3k�0*�cO�����5ne8T(��vٕ��S,�Y��L5���%��v����VֿV(r\_W��_�W lX�l[�NՓ�����Bb��	���0�؄�r��Ti8C�r�N��{OK̄O;�f�z��t^���6�	/n�"c���unNK����;�W�M:��In���z2�����m�	'J"t�Wd*	j8��_9�X��l���,SY���Y��P�2��M��7���� h��-�\Ϙ�m+.$ݭ "��࿋����p�-L�ɮJ�py���wn�v���#k>�����(ט2�^�rb[}"0�A� #+�:g��:�(�K�w�U�$@չ��NQ�n�^)/�hB��=��J�{R��E�N���8����zX�]��6i�#f��T-�Ŭ���zϦ����S�e�K���+�2����� ��Z/�-]t��{��=,t��6���9���@׵UЙ��+C2��h�:Y���)Sj�>W�v�c3��¤�O0�+�u�BǴ!�o���C�~���X����Jcenq�BGE"H�7-�Lt$\�s�T��s�j�[1�5>3�W�ND��J#G�k������n�� �����Z^69T��Ć���Y�a��U��h^���a�,]�������i���c��2ƽ�ԓL��n�m����1�V��3�m+�̭WyW�^�=��"$fB�3�ʏ�L�Jc��y^�� �Y[�R^7?�r얝�*56e<5�F�A�e��a�}���Ë0&�4�J���}�gf؅��@���+P�h�Йy����r���b��Z��S�<���7��v)���̳�����W�{H[�V~�_���D٥t�J�M�{lQ��%��IY�����B�Hd��4���4��=�ϥ0����?QOC)����f��a"1<(�2x���T4b�a� ����CP��zRY @g�x��`BV��X�y�i'�;�Jwr՜���}_c�5��0*%MX l�� ����cu�c�uPW�� ���*����w��t?��3@X;�m�g��^�`�hNc�Q\������ΰ�pt4��ݜ}^ћ�^Y�P�P���(��I� g�vĬ����gPQ��7G���%�99A]� Bl�H�ʫ?ϣ2�n`d;�}��E���S��� �4�eo}�!��^
��,�L5G���݈6��:&'�"�&�'
|j��]BeA�����g��H��3�žm'�H�Z��7��t(�;�c'�(�4�Y����%��:P.7�օ!�ݟta�����g>Rq*�i������	ѭ�5��6���)1�1��-�▆d/�mق��x��yW�!�9�Z��y���K���hr�hY�^��.�P���,�S�`q�
e�jG���"^���*s��cP�����2��u-hxcm�q��]f)�}l����(M���ծ�t��)P�p���8ff�r ����v
G��������f�ò��3��f�ժ��
���(�]�w�
-��)R,��ޒt�t$�%u�@�:{�KI��a��LŢ�+�5�&&j��c�Q��֜|e���p���#��'dS�Ie�x��	[  ]o�ˇ�E���).��A=5�/����.Q?��X%��V�M�dNA�{e}�k�xQ�K��Fwbp��.Pw��t6��0D�`�K����j&�|CEŚx��1�!jY:C���Q�Y�;������|So��?sXo/*QpϚ�Ԗn�?>Ya��f��@��@w��x�<]9-N!C5��Z�_*�D�a�;�]}2
̨
m�.^�z𠻚��5�Gm����!}���N�g�Č`ط�Q�� �_�!���F��6�(.ߑv����_.�C^�uk+�x>!:B�8�G���oEC��y)�>\�H��_T���Ā�D?��`��bRM�3*=�:6�ى�(9��\��I�t�*O�|'��9a��&��7|&�V͡8a>J�u�P��2(��aJ���@xF{�Q9���1B��Ҟ��}�C�sh3���F 7�&�^�߱��]F�j�Z&�)l:_�Ӳ��Iؐ&�)'s����|����m]�;�D^OQ³K\�!	6}i�TyŚ�Whd�ۨ����^��B�o��B�R�tKW���~�<$�Ȯ�V��[HA����Y(a7�~R~�|���j���TR���j�����o�ۢ��ro*������Xf?F��1���_�9A�"�U�r�A*5��I��1yl	��	i%b�c�.�H ���3�͐�={v����$+�f�,aUN~"w���5�1Ѱ!
����A��ܶ�.�6F޳�a����_��	D��U�~�%T�e��P֡�/C��Ai�y���;SL-���A�z���Z��&��|�K��)�ݚf�p'�������͎��}��:R��������.���\��D�#��
C�����2"=�<�h���UG�^��_�܍��}�:9m�ao�ML���fͺix�$a����C�����@�zW��E�����WT���¤�)~WyӅWa�G�Ǩ�sݡ(�����acP$x�/��"(�O���J%6�p��0�o�����<��ұ�� �����	GVq���V�^`{A1�'M9RLC�°�=k�ٟ�IP�x���k�t�U�[�q��Kn-�Y��{��5�Tڈ?Y���.��6�r1عg���|��E7�e����1V�h8�4��,ö"�NQ��"�^���=u�v�:p�H���o�Nz� {���k�~
;�:#N��p�i`�>@����E��YCs��cMn��'�O�T4}C�����҃��S��݀��~3��I��h��������y�P[���~�-�*��L;l�Ec�uB	r\�-`��������˨Y��Z6���7�7\����C?���/��ڜ��a�R��,L�8z]��m�34�w1���Ӏ`|wvo�G�ǉ�R����A��	��4���7�kV�=ʗ�]�A�Q:��cK~�	t���tS� ���v�0�^Z�6�j ���Dg��L
�SdK���R�(�>� 7�����h����L�"7�.飆Uٗ�PΕk�*��#y=�x���,=�sZa������j��y�������%a����&���)�djg���% ua��AA{sz�5Of���QT�BBo�ޏ�\�#��hqN��:��vN��ǒ;�˭��O��/_�2u��|�d�h#�Xg�,/�����Rg�k��I��>eS��!/Yv��|y���,y�jKG+u����������"����VF0�"CzV^e�hh�a��K��ݿ�3G��%��į�׮-D
�����_�j��E�{2V�iэBJ����0oS�x�Z/G�k��9D��O��a�&}x�"P	��L�I�1��t�R�q�j�!�,_d�7���3A���%����*~���o�8h��u����;�e�W@�A�������"	�e��'�T�rsh���(�;����p|�IA�� ��̷��9�5��im���X�o��]�0,,Y����/�B$�����%1���9<��'�8���&�=P�*���B`|j�iL|�mNU<!F�	t�6	�W����_ɟ";�ˉ�*��4�������R�@x�=�qɋze��ռM��9!=	ߕG�ѱ�C=g�����5~�z�e����~5�b����OJ��|�S�"�S���r�?g���L�q�Z��۴�ܨ�@S���0Z�L��tF�P���lx ��7�%�|"��D���S�\�pzlf��8�{��Zv��=��8V1oU�0��F�A�c Y{��'2bC�W����}�F\��&�3Zu���9CË@�g�z��:�Z* ��w��o)��5�Hx;6n�W�{�y��:��v����;���C�G4�N�4��g7y��c�a�l�P3� ��8�vFl�nJ7_�|��U�(���|x�[~�Lci�z�eƳ�˕5��~�V��]Zu����o�"�	tR���Y��a�G�4 |՚P�V>F���j�rrK&�
��+����e�,ƧG8��L�}��܋�c�*���'K؁?��>��S7>8K�۫�;��쒁�ߵ �����`w0�_���J�	u؋^l�G�x���Z[hPd��R�L�}_�p��ǒ�pbm�k�Wn����zWa�)'�:��2��*A1��q<��2 W�Я�Ѿ^Ш�ꅅ��u�.?�
*�������8i��^4+�L���?'�Љ|C�T%\�W&q�ˀ���y���(/�_�����VlC^U��M�=�͠�n��g��%�WEr�v�&MQ��@��0�H����A	sT�h��F�~֦��cv����'��ql�]��C,�qȃ�))�ws���} v���U��ϟ���g�����/+#([��j0uT��{�jD��Qka�*.�	Jt��E��y�|�fϺ��#�2f9������PZ�Ci��B����@9j�Q�)�t���\�C����V�~�,�/CSN���(�\�X�5]JuU/�'�\��~���]�A��v/�
��
��2W��Q�B�4��jJ�����ꬉ��Z��O����0ox����՟��v��<�����"��0X� ~����{ܰj��A��#�o��2�@�pL0N��6������)�c���C*f�el�����M!�PT�4xΝ�7��#ڔY��:�z�FE��z=������$)��!�-�6d����JM����I�~^g@����Ԯ�.���M����pÛߞ䌥�3SV���9����n������;/�n�`�^kSqg����0V��5#����
Z�L��:��C�]&t�������I̃Mnq�����k! �'�򳄸'?s����7�F�8�m��TqR$uΐ���O=��u��~xC�_̸D�����i�nE��Y��n4�*��qHg !Dm�n��ILN=S�X ����mB�N��B������U6�i	FS�1@�1���D�j���ׇr�[�NL�W������0%8�Z9.�#��G�B�+����(� |f�u����56�^X��ί%R��Cd�Ԙ*��,K��K��d��-�����ЀcڐI����L�)��+��QA婘��ٿ�UgK�V�4� �>����h�O�p9�|�L	�Ȧ��f��M�"�.�B��L�b��>F?�.�.h��7�6@S~��&���m:E�9T�(R4��AM�p�`b^S�*�v{I�?�U$]5�4���O|I��p��4|�^Y�/���*p��ε��3���BU6Ȑ*����F��T�����ze
&Q�6b߷�Qm����(��x�9���0���E���I��6F����%jfr��!sM��xr/�I)u��{�Th5 ���e�R;%\���t5�؈S=e���)NC�a��XѬe����b�*$]�B�A�8��2S.v�6qF�����,z0Z��F�b�'�@�`ڢ��L���	�l�6���tИ�N#T����z2Ojx4�?����p����E����'�7�,��C]��I��;ş%we�zUې��^a��)�e�>_�IyiSv�RpY����)#kd�}QX���	���F�S�b�P�#|%�9@m��2�j}i��n���2�5*�Q����|-�$��vj�i�F���W�$�
���x�שP��P���㾵��S���`2z�!�h�I�*�r+��2����N��e39�f�|jj�,V��q�� s�k(����BUGs���lU@g�����9�1�z/�dW��
0�-�GX�Phh} r��߂��D|ዡ/��JDX�\l�%�+j��)�F^M����W%������$Zt׳�׉��c����/�k_~2J�,�23l�$�_?�W-�/XAn#��Bą��&�k<z�EӁ���mX�voR�����W�f�����Q��Z�Os�vU���0�*���y�_졪�{������;Ԛ��|!�[j���"�S�5�����2� �/hV������6��	&0x�McPK����jh�az�7�#��.!.�]Ⱦt�h"��7^�W�l����Կ?^�I���y��q�U$�.'Il��%U6 �X��(A�B9�I���~q3�m��}kr->]��)4�ބ���[ӏ$5�e��>:BA|9葅�+/�[��J��n�{���r�YW�1\G���F~eW��4ٶTh�� h^^�?6�mس��E���u��dw�9��H���-��.�0�iEϾ�m=�}}��E��ϮUW�)L��5��`/���}����`���mRN�m�R�\���Y�#�����g�V;��a������M��[��*^�%.�l '&�0T6;�3�>`�8p�Iz�	���)o#�/�Pn��o;n�ibI|-oi��kOޕ����:jiо�,��>��[up��=Մ�Zq�DB�p��^Y� UR
հ�"i���Z�&��J׾c��5���`ru\��8zs=�j�~���k8��q�����HN�h�
:_G$K���6�|Z��(0�i�;���47dpd�W*cмO);���/z|�˼R�h��#>�+3ω->>BڸB5�����5�C�&�p�,��H(>��bs�mTW�YY���؅�LsnT��[y�Z	�ױ�~��� dj
��)����T��hW]\
P�쌌z���V�ׁ��8����y:�f-ܹ��`p�!?o4)�/s�r<�rf,�Fu�;I�(�����~�Ń1N=U�g����Ս`�/��+�W2�`�yR2nt��fN΀;GɊ悩?tUL_[�!��ݕ!?K�:L	ӳ0�CSCe(���Og��� ���u���!�aWd�����1�(I��S���g"��Q�odb��А�Zvv�c��Q*��A 1�� ����q��~��pa�ұ��8��m(.�>�C�# �O�9�;c��n��A�w<�C�'�_g�X�~��t�7KWW �ǣ�@���� �@�������EL�%L?�}���3����AVp�b�}*�=�D�sHװ23F��b���R�_�'��I�r��&B�Ñ��ڨ���7#�ڳ��w�Pu�4Ǝ�utaT7��v#�R�Zn�ܯ)f��Mџ��C�jZy�V5$���J��}���1�A/�wJp<����	9��'�$_�2��e��lߣ�@��&��B�<%�����f�q�GIl�9�Ǔ�&����%����-]-U�;��*�=-�_��0��-)�S7�e���V�F۬8���V`��}uIz�;)R8������;���VR>���3�2Ս��Y��p���z�"���+��,�a��X�o�6N�[T������ר�;�2��C{ڒ0�,�DM(�9�Z钊H܉5h�(��/e+
�Q��ĸ~w���j��	��|��}%fa/�c�H�A�/j�f�X:����<��)uQp�O�.W�>���h�M��.v�aO\!��=��ݽX@s��ʒ��O��'�����I��F�9-Ƕr��}��T�)��ք��m)n� R�<O<.�@���GNE�:��SN,S��^|)�i��<O(�8\C��N1oY�MU��0G��M����5��y]�$g9M�7�P-�v�AA���Ե���y�d�BǼ�0�����Vz�%bΣ�'�V��K�Y$C���e*~�Ne���Y8+�r�1/l�1��jQ4��Zw�5����
�x����o���&Ń�@g�Pm�+G�xV'�6vD��S��~�z,�Sќe���
W{D�QJ���3�y�ow��zD�ѷ����v?��	��� S�����9�t!��;c���D	І���1v\ڵ��N�B��fEIj������ajŒ��"K� v��e��k�J���l`.�@� 	0�(Iwv^d*�b*�u�x�z�3�@q&(��7��n:U���?��T�!�rA����G�R�̦�SNV'�ҙ���2g�4���؍5���o�I�+>���6O)L_+�UE��
DY��<�w�o+������,"�=E �G�4�?W�Hz��@�K�'�Kzf&
��M�}IJizÆ�E�K:�$+Oqx	,��ʊ����35��E�Ε�B�����Z�V�M�}.mͳً��噉F�̙=���]"WQi!Br���{cLmݻG�<aa�,�ʐQM����	��T1'
�u��r�e�+���cE����̈́�w"��6�&�'b���k�Y��2[����>�1�0�����Ǟ�|����x <�[�o�(�;�؁���p>�9#��~w�!A��|,���L�Qv"�V0�U�֓pu6C�I�DD�-	B�-I�h8+�'{�E���Q
N���b�Kw�}�&u^�dz��	}�+��z־�=K	N���h�^�Na�������I�MZ>t�#'a5�1� �Wt�O�=��S�!�įދ'2�ܲPȕh�t!;ۯW�/�Ō=���e��}'n>2a��/7k����1yga\� JL��1�wz��]�s>lvuņ;d
�t}���s�ԗgy�����w�\yeӦ 4�R�00N]$P[�2����xt09IW,� �`�WᲙ_� 0m�������S���Q�ް�Q�:V�H3���φ���5��,%�h�98��B�RT�W'%x��v?2H�>N�#�)� ͘�*ŸE[��)�4m`�Yvt��GDf�i��E����F��*Иá�v�j�7?}󨫢��Ӕ=)�n.��P��{ ,�hL���0W���U���(.�Q�WU�Q��wk!<ݗ«Dӏ��ͩހ�BW��kVLcN|o�{�Ƭ�;k�B:O%����`��xū`���s��M@
�s=�D�&��H�f�Z��20r��u�P�?����F���&�ނ��y�/C�$��ӽ�%���7��9U�$d3�2����E���	��_�ϓ̫�P���Be%y1=���J8�Gǳ2�s#��� ���zW�yi?l�c
ҷ�F��A����"[�Ex�
e�r{�X2p�C�,���~��E�~���#�ӽ��^<�I�1��e��������߽�l�z����J�4�W����/�]����c<�ſ����Q<G����|��U>��h�Qk]�_2�b��iEb�x6�s�c�p�Tm�6�3Y��r���Ѕ�E��y3���+���r�jI'���M���\02���wfh��Sߟ��b%��u�F���s���U����'E˓U����O�t�|܆P'�E���b����N~���	����I2��2Y��L�d��?�J!�Ͳ �(�� �>FV*��Pt�H����X�h�l��lt+��Ո�{qiosa{$%d�� ��v:+[�&>	�=B�gvD���i_f�F��P��I =Ә�ŵ����dc�{���Pu�"������Vlb<c�R*P���w��G�=��s>!��$�������3_	c�4�B��.i��H����F�^l�>.�&et�#6A]�ޣ�W{�E���t�]�c�.��I0���)�3��F��~��C�!x�?���N����T�3_?��y{#���߁�&���֜ADq� DS3"��_G�p)�J0�P�ց��d�Y֗y�J�_1Ӣm�Nt����S b+׋Rxݦ'�#�/|��9B"Ɏ��0��+W2�
�����t��y��l��'+-EN��U���?SX��}�=�N/B�����tYP
�7C�g*�'��2�<��W�8!.����a�3�ܼ��R�n��/g/��Q����f���X��!,ޘ����P2�K}�f��>��S��f�[��apYB	�^VʫCWDc�gEbW���B��޾F�Վmr�1"���Hݩn�R}W.y�H[��<[�`�9�(�ޭ�����]��G̖��>ȵb��W�l�T_�^�ө�N�c}�!��t�RQ���q�B.P��4
fyd������_�V�܂\�8b�*� �T�J�t�C��|��Y��b�(��+0���v�8����}����Gu���Ǡ�~8�MC�>uc ̒N�|�Ƈ�{1X�[�%��޶5g H��r K��_���g?Wѐo*�|*/e)���Z|�)��d�sp�˦�F x��O��W?���?N��j����\�MvD�*]�����d��NE/�y�US������4�a��Gk��u�@����R?�ta�;���)˶.�K�L5����7e���;>.��[^�~���0%���e�l�W��-�S��x��=,`=����5��&Prl�+H��p�?#�la�L�i����mϞI�[[)Kx��vf�A�+aU
e8C��KE3��t��] ��xs��:��Ӿ#�H�� #G�a,�K���)�(8J@���c�
����պc�%��*ġ��� b� &�^;���3�H����8ZJ<|!�ST ~]pߓ��z� ���EF1���m�l�����rg�?*��d�������Kˑ^m�%Ұ�=!�VVW̵���>����6g�\���=��>7s��rt��T��R2��~�h���G�kXs)s)��EY�\��^^+�H�>��=���D�����]#�ƃ&��,d�aPw��6��z���4�?��URDbI}�Ӯ��Ϻ��N�DQr��\0�a�[�MG�Z����P����?�*<B�����9��q�#�lNX-����Qֆ�H�(���4[������ȲI�1�ʩ��9૨c�ߛ����گ�-����b�lY��_�gUg��������n���{n����n��x�IO\m��t���
[�0���Q��
��U�%jM��`xG���Ie)������� ���n_EaK��Z�U�?�F�v$Z;(W��T֩@�-�|{�$��4o+�:��F����ϻ�*hX'��f�ǆ�XMz���]��КE=zB�����E�h���X��s��Z�m��;�`�*�����ɥ�u$eS(`ٵ|J�̄��D��D^�U%��$Wc%v���Z�kw��N�Ԣh��\���F�����Q�Qk%��)��Nߠ%%d�?P������3�����)�������oC����l�qvQ��+�wWF���齱��w@$�����p��'����\ß#Q�э��J�p�I_-�21����J�$<���r7'Ơ��Q�E��� =5#�r�5HS㹸��BJ�8�����#][�����v��r �|�L�0H�
����L�x�m��������_nL���0�n[�����d����/���J`�JX��Y`��@
De�ɬRa��[��̚��U`#�5��׸D!������$:"K�z�W@����u�`T@�!o$+���P�OAp �{����/n��%(�i�
g�⺳�h��)�:>���p���/7��}K�����|��[�����-��j˟Є��d�4��+�r�qHR�ce������{ؼ�G�%5��y�%�$<G�Cgd���]�_��G#X�L[MS��ijn����̢�ħ�]%�z�S�D/��A��P��Et]��F��[k�`$�+�$��$i?|=��$�l�)T2
b���h_ 5��=>��7�/`"�ހ\ۦy�^�5<�0�\X����qε!~U�ՙ�����!ooO+��(��&��Y����eK�}T�:a����R���f���M���h��e�Б�~�U��;��IX�+��͕��%AO��Sd,K�4�+��B�3 �f�s����a2�+]�C=� 3aJ��(�|����4�n���K��ʹRij'�Ri;z��Ǽul-��b� ���6cm�?&W�%1T&�# ��^��Rhy�L��������}H��V�'G���1TȌIM=��a��ȏ�[�(���Fw�i�u ]�6�,C���i�J��W^�W-���p�k��bf2B�f�N�RQ�e��l�z��ya|HêW�H[f+�d%�1�c�DS3�}��
n)e��|yy�\�%Ik5�>_�`_ZYy�x\��� ��lı+)��Z�6$B����YC�rdh��rm����) �a���?�#8���!�5�<�;��C+᯷���?Φ�Q��}�B�^)l�2SA�6�𽔾��Q��ς�/�7��٪���[�i2�6�,
��dp�_�o&r����%e�4�A}~��N�(\��b��P׼ڈf����R�*&��%N`q�,��S�L��-���r_��+iC�^A�:@�j:�Z��:�G��ӿqthq�B��N@�hq�V��t��c�xv>����;x��}��?�) 3<&�i����A�0������W�ɲ3i��>��yH#���|N�S ����H���c�e5T�*����&��'b`[Į\���exۃ�V�`$$����6���/����C@�e�Āӝ#���DJ�#��
f�YIH(�$�@I����Р��������������.�_et7�8���@�B$��ǝ�I������<@J���@*FO��>u�׏�7��ٕ��h���Q��Q�^x��A�g83P�v��r�qm�lQ��'����	���^k��S)�UP�H[��}�%j�^��%�� ؠ�0�n�5����!�F��7m�Hd&,Ow�P�ǝW�C(���������(��m��OnA/���ϻ>�RU^繢���q��G���6�?; ����D�f=�=�A�X�}�z�Yo���j�8�0��t���gH�|<�}J�LAt�$��qu����R2JݏZ�H!i҇�~��xu�65!��]��"Wh�4N���д�b$+Lj}���˲[P��$�ҵ-Kϫ���v�<7�iX�՝�y���@ PX� ��a�t�~8y��pK�:=~Q����(c�!���E+)N�����ȇ�K�C˰�Ym�Y1�ly}�-�ǦSpU�ݯ��~m�k���ĵ���U�E�@͙6]��tGJL`R��S�%��q�1Ur}�*=��Z���5�d��.�J�@T�vvb�v�z�&Ɠ��j�g *�����H����*��N��,���F�o^�� onf�*��Qdq���AplDCX���q��L`ɥ��6d��rs�&Xr��*/� ��V���>�>I.���泼aEo�6�0�ކޡ~/.�%��N(���zBi=�jg���h@�?r��N�P��9�퐲߉N�]�E���p�O�N�cz�;������Z��ԊZ7�i��Ht@o
�6��]2�׫O/�0�����;-!	�>�T���?z���5��+���T�b�
��R�<:�L��k;5�T�fSt��Ҷ�D9/��&�k�5�5(��"����j-�{��jJ(�y�*2kH���n�V=��7Jе����/b��#����a<�N�rK������V�0� ���X���^��ȷ��ݗ��0ݛRCh����rڭ{?+"D&p$��%)G�(�_��p��!m�ѧ�!����޼`P{��LG��U@��H�<��o�H�x}ĻK��s�{�B¸E2&J���o�A'� (��/�t��2Mq�cF�a����\^�y��J8v��6����"��ns�f|Ki������Hq�d��M'O��U���~͔�$ ��zS����9d�w�&1��~^P*�)8@��]��2��ĭ��Ȃ�����3E;{��ѽ+2����I���|f��vt�K�'�-#�j:;>���T~<�O�ဵq�M�TzN��J��	�������U��m��i�zk�FTF�K+�M���f��h/ڈ���M!Iе�L�D�q�Z���r�M���RX������Ct/<)��8�����hA��V��W�8-M��(g�o�KRٖ`G��q������<,P��7�|�y�"P� u�U�B�%����O�"�qD�3��0��J0��(��_Գ�d��AZ	��G��GOq����!��V��aEk��T�@ɧ5��E�z����썞�B\*4i����^S  �Mc��d�f9�^>���$��2�p�i�݂c�BX)�wI�C_kL �=�v�i�>�M�wQ��x�^�5�S��hu�n��0[�8���}�&�0{'���p��N�!T�pB��"�F�������%�$�4�jJ6��`�e�5�kW��>`	�Z]1`K	���ɟ�HkO9k\gT�n���KL��S��z��{��sx�����*���X�_o�����A����KW�|�>����0*�c`�z�1��,�n �(y����G6� ���Cy�mS�S��C���Q��BEg�n�ё@����Scw4^�2�@�*�ٍ�_�ap����m�m�2�����P�M�f����3��� 3��B��!Aϱ�o�I��2�-�*ԫ���d�������Ru�;�է^��9��Z�dP���7F�)k%����Q�y���<�N���Ef�,ԫ����۶�>8��Z[���P�X;��ŵ��{@�])��	�%�=wA�g���刐G�H�!��yc����|$l�E����D_�&AahŔX|E	���gaCUf�~+�L��C�ݶ4!�̋��X�1'f�+x�Jcu�x�ˠc!E�&��Ix����p	����}u�О!XZ	�3�*�tU,�O+��q;Ҩ�"ˣ��ҋ��p�3]��t�9��zL�܀<gy8��㸰����Sxs̻�'�V8�մ|�/�KrK���!
��t��9�pe@E}�m���>"aa�A�Bi}�@^�\�0E���`@eFڧ����X���� Ip9��R�Ȩ$�ڜ1�R��-�0�d�IX���� O�����B�:�v�6���L^E�N�}*��:x[��>�����5-��a�,l��4&�x	���9�5��2��crl��G>�$5��L�
���B�Or��A�=*C�K���j�A	��"IT3�=W����Ɋ%v��Am���Nð?�����~�^�o�glL�/)4�%Xo��cb/K(�-�_|k����[W�+������~��/ϭ��5&���ѣPY6gHm�j#V:�h�9��>���U,�E8 �İݪ�ee����(���A�V�h��mpR�C
��}�6���ܥXo���; �x��h*_�����k�߯a��r:��G�@���k��7=NhV'>U��L��K�|K�*ݶa�D���'#N�\!-D�q.��e���u��S �����2��X8�G2i�0/��CЮ�h�p@{�q$<��c�Q��&�u�ǡ�xH�D�����i�����f����"��>�0_N`����D��?����둼�r!����9;�#�: �(���ˡ�`��@[	������j�
������m��� ���mʙ1�<�+�Ҙ�v�߲��vm�k��&�q�0+sB�
d�V�Y�ɂG+�Mj��=���Ӂ��a���م��( �e%	)��N[J;��IA�{�Q�c3?M��80P����؂�ȹۼ`a�"� �Q��i �~�u�:Wr�4��J���!z��udq_}��yn˷�J�_x_F�_�A�u[��\�����M�˖ ��P�#�"�����K�9�ȇW.�ݴ��r"�	C���y���8d#�ʎ��۴�F�EC�B[��<�����9�%߸ٓ2�DuT�����+��q�G,����h;C��B�Q�/_��բ��f� gf*�}��o�ƥM��cA��nW��+VO���$}����ix��V����C��b��&Lr|��Y8m.�2hs"���Th�8.e������f���X�s�?S+�(j]�o]|�g����r���ǰe�J6�y���)s�e����M��H"nV�w���ѭ���AO^
��}"/U~����������9���oKh,�ƷA�ZR8�]� �p��f�s�Ǔ�}�<Y��%��QL�k������.bl/��.���D`�N�C.��1C�iÃ��p��^-��k{&1�1��%�Ċ@�	ؒ� 4$o���|Ľ5nv\3`v՚�,���߽k�X�hEQwEJa`���;���G�w���i"2U��g'�$��"yFd-�j�]��C#'~��92a�� F�1�ꍉ�h-�ˤ�l@�I	'OK�ȳ!�|��c�l|�Gdmg^0���X��_�Z��T�7C�/�b	�ب����?����f�����6��AJ�K
Mގ��T9^�W�f3&��
�q]�F�*�s���\+ژ�G��[~���+����H��q��^�a��Fqw����� �O���N�Qj}�M�r1@}�G�)��}r4W=�[Ok�!.���q]���)q��<����쀠hLObHCUeXF+	���ӹ�hڶ� �.�u�E�m�2?��?����A>�+��%T9 S�ܔ�"}�w���L&���R�Bd �F|U6�UWα��#�ՠiÏJ�*�
������H�4w�W됯(W����X����"�$0)�"WK�.�,.y-�ϊZW%	��e;&���]��|J����ū�o4<�]�1L	�b�3ރ���P�-g˃Nb�k�hM!����JqJ��l5���W���?h��i�ӟ��u�y	�a�&U��&��rřpۡ?�:z3���S&�[׋�-u�7���,���8���T�ʄ9� Uf��X>�\W�~�Pr�|�V�~�;���W���q�9�K�<�F��əqBQ�4��`4�;��U��֥��&�D�U*��U�|�w1ቂ�xG���Տ�.�|¥ݍ��h�E1G��LӞ���8�R��B�e夿Pd��V�;�4���#�kK�"��y���%1�BI���DV��o�p?b�0M���?��� ���!�� I}#1'T~��t�6��.|®')����ș�	d1����0y�eR�p���R�~�:�A�F����>ɷ�~D���z���(-�ǝ�^NZ���p��m!�PQ|�jXΙL��~��n����1׆ztU]��l�T&��l1�G�P�֦�ڌ,Dq�֗�h���0~���*4��:�Um�ۗ4(jE�r=D�	�:Ǹ�h����/aZ5�Fo�	m@%�^��7�ƛ�6W�o!�p���Uy�E�Z�#h�����ғ�C��_��B.���[�P:O;��C�B��p�+���\��u���qW�Y��N�~`ғR�a��q$�̛� �H�h�6�xddp)��8Q�`�$�B��7�*��+�N�8ÙVŠh���֘;5�����G���9!N�I}�|�	D�u������f�1)���:#��"I��:".j��I"O?�1%Œp'�2��̍-�rg���ү�(��3���?CW/v��B��FH�˱�"p��\pv��z�フ�ld�`��bf2���F����x��3�垙c��*����{:�.t?����lT��E�Y�nڣ��$}�&ÖY6�Z��*��ڪ�� X�T5F�:� ���z�Oy���U�k>tiǳW-\{1_���i<H�rw�*��lL��7Z�Q�2pHɱ��m��8QYR4ͩ6�/�q�9)OЀ��x��(���v��%H��TfD鉴Tn`�w&�b������������ZR4j�#�O&D�j+�G�N�����yN�N�@|��Z��5��d���ޅ��U����N2�nf"���]�����HA��A��|�p�F=\��o���G�לK��9��6?�܄�n�>��g1E�✯��e��n��Gp��>/����ϕԌ���er��GCJFǤ~����E��8?�J���ܼ���i.g/TC��ٽ
�)a���Z3��Y�I���C�ޫ�=8b~�D>�$�U����l����Qfz$R^O�-g�qH�'l4��n*�^;�ܗ/z�W$�V_b�Ro�l9P#��R���[�q��7ֹ���XVQĴB�do�}S�X,�:;%�)��μ+U��kow4?D���_7�9�*0��4q�$�������M6�M�1��m\n�wڄ�Ӎ�}匳x2���hL�%��N�u~$&y݌"=�|w�,��;��Z�C�(~8Q�z�����x[�*c�K0���3l�6�e-��{�M����A�qm��ǳɽ	ֶm�y�-�����`��LV���k���d^�f���� nÂAp Eu�'T�����	���?=7��Yk�k�h���Лᒀ�k{�}��O �6��8�'w.�5�۳�U��9a�bv���H�j��nE��qܗ���'�?k�;#Tm�Y��c���>R�fյ&��d�lEk���`��d�t�X���*Q���������T�c
\���~C�*)�~���d��Fы��\!ܭ�(�=5��υ�^�GI�GT=zr�Z�&X9�$�@ȪO��G������{����*��	����$,���&�*\�[t:y���hwbG�su�.�ɝ
��^r�Y���f�l���@���a��BR�U�<����8�)�����e'�򣦗�T�����7]K��<��Z����Bꐐ�	��{���$Rie�yYƟ�JMY�1�	
ߦh��}�x��l�n�ڕ���[}�&��@����
�Po;��Gw����L+�&)Ll��;w?}o� �/\�Jm@��"9�a��;Dw����]������)Ӷ���;x�����|�,�O侤6$RZ캼c7��k"��Ӊ1&��,+�!�h�ɯM�[U�9��������e�c��1ɗE.�\U�i;pB�e�نө?�n����Xd_DV����ڑ�R� �t?��<��tY5<9�='�*�)�|��e��"��7��4︆�C"�S��a��z
e�-��0I�{H��I�9��w�˔϶m��=��K�ৎ.�� �w$��M>ЉC�T���P�b|{_��hm�6(οۓ���<�`����۩�7����ǺH�X�ʳ��_��G?�<g3�����j��kO�u��0j���d�ĝ��~��	�	~�T±�Y �w�~�R`x�q����N�qa$�Mp���.��V���OZ�L�yZ�E\.�mf-�8�0��Lt�k{��O
�΢~(���PT��:�~Rf��U)?�F����yx�[���8��_�i��T�2ٻ�����ŭ#�c��G�T�*O�+Ln`$�K�Ǣ�"��,�pC!]=;�9���V'��$Gٴ�{�v�&�7�Nd�֍�;Ω��Ֆ�2`9%���N��^�,�e�,pnzf�^����^�����\��z$���c�M�ǳ@7/>ɩ�k��N0� �Is�BƸ.h׎fZ�.A ����G3��Uz씏���n[+W�a짤�ҦOn�]lc���b$�5U��:��r�K=2rp�α��1v����l�l�B+1!�; �����p�������}ퟍ8�<Ծ�]
K���P�m�Fz!}���}���k1� nG���-�0&!VctX�#@�7U<㍱��37�P��\r�^��MMR���e2��$`��ҷ,B��:�۝Z[P}���5��'
�r�
�w*m���6���S��O�70B��d�
$T������w��_���6&iB=���Gw���2�2�pc�q��[�ڂ����U�O���D�)�q��n�X���x3�/�m$]�Q�Ӝ�z9�[|h����	��8d�
�v6<Xކ]�����A�v��f5��U-��s�h4��P��d	�h�64E��EY�C�$��`���(/����:Ǽ��'~�v��e��9*=1H1�855=�b��j���:Ji��Q2 u�AR�f}���������5���xPכ=�vp��e��3�=����^�!)jO��qq��2���u{�G��x�x�N}jy��ܰm�͈:&	�. �?��T
���\�Z$a����Y��ֱz�g����X� �6�U���.�Ma����|�#��(���i����t}�Dc�] =����{.]	�~�s:5;v��%��X�jcΨ46��s�.A]!x��/7ίc�y|�7��@[����D�-�d(.���|k��~���[���f����Z%���}�,YO��*L�ťf�Vym�5�{k����:���o-��$���#���3�!���0�W��K�Ŕ,�3v'�.�f��� LbI��}m�u3YG�r_I�g�GS,X���ڢɤ����5`͚�����x�[�sx�$3V�*1����*Z�W ���li�ʄ#�%��'0�iͫɩc��B�f;�޻̯|M�^�:Jm�
�3���O��p�ُW��[r3:�ϖ�r?r�KC�?8���w�.GNA��i&�{j�W<(�@ŭjB�K ��pH.���ѫ[�:�˓�c5�z�*�b����=S����4sc��&���5��w��Գ�@���M�|%D@�nմM'pu1�p�s��>���T�G�,�@@0��2u�:,!����	�r������ Y��j�������|���oO���'h�����"u�/�t�u�b<1���
tȬ�D��]F�[7��W){cR`Z��ԣ�'��ٝ�%Lg�T*�j�/j��������]����������Ԣ"�E���tXC�q~�3⃒��:w�JV̛�\G4O�k���e�����?�lj'n*Z�@X&�|tL���:��<�V�P�B�M����-��ZI<��J\���Yєh��`<�b������%߮kwN��'7�#g��"�d)s9[�v��a���2��Os�]YT@�渝8��r�2�c�c!f-��*az���m�uF�p;	7×�O�.k���ɟ���@�K2��;���=�4h-��^�.໋DU�ƴ/����!�T�E����l�V�]都�h��x��9�9'��)V�Vb�A�m���6Lx-N �Y��χ������0���e�Ԣ,s���Ֆ
.���򶤰�����P�
�ҩ����9%;�
���������!��k�Jv�G�y>�J���2G��7�P��+�p� �����or�����C�W��+V]�#�N�l�O����6́�U5?z5�`�V^Z}$�Q����ʇ;�4�Ի�������}��Q���&��-��jɝ���WNܑaWQ˷M��1U�K��Z�q��m�����c0��Cy��t�g�`2~2�Ŀ�"_Mo�K�k������LXk�ޚw1n$j��n�R$�	��%�F������L���ȳ2�5�n� m�����O6�&��4���*4Oǳ	!�Ł�mX}�-e������C�#�`޾{�}��
�1��I,(�

���B��a���5��35c�Q�ѝ���o7o܋.f��43��c��}�L O$Y������p���e�s�c�3n�����W&�/dtw9�wU$jX#/���N4o}}=�f��vv� ���P�iy;Ӭ3��س��U(��BKG�vڮ��olBJ��%WL�,��1p���T�$�[�.�ܢ'���o�`���5RP(�qX�ۈ��9_�5Tf��p��!i��sC	aI���Wa�<�J�wd0�����{G��p�9��H���8�tƪ�s��$��0˲ �~rfz�^�(������t��Q�X���{�X�/��p���yv��-�^$cn��EC/��m� �v�Dd/��=G74b��Cÿ0��gm�SK��g%�����Ԥ��o�������7�3���z��T�2�
`[oX@J�<0��ܩĦ����%�.5E�z3��;J:m�X�`���O�|D["x�՜히Ą(���ɩ��f��ٽ�;���F�̈́שUA��(� �I..� �,��J}6e���B�ͦ��?>����B�sC?J@}	��b����!��O����a#>ٚ��. :���L�6��"k���6.]��=A!u:Z;Ke9Z���z��5k��˝���m~	5Ǹ�X����)t�wѳ���H"y0b�+�:�� �u�����$��ջ8�SJ%F�l�xˉr�9�J#1ݨ���󧔃
(�%���}�| �C���8�%�Cj����?z� ƭ�y��3��i�V��M��t��e�k����k�iC�TE�D�e�/��(����v�d�M+���Ԧ;���AP�;l<�������C5~�%ٮ�Ju
���Y����&�5�鱇�G�A#��	I����N���G��5����?=+��a���o2�c���vP}"������.��~ L�ud9X��t��%�&��K�+��-�pG`��뗱�1EW��#��ƀǊ��� 7)�Po{]C��`h��O��/���kI=�@���P��#�o�,jڝ�S�A^œ]J�m���dd[
�9"�Ϧ��93k�5O:��5:S�4��T�2=���~t���s�G��pC���괅n+��qdS��v�`O�l���	��r��-��I�ŋ��T8e�)q�p�0���YK�� ���ޱ����r#�(ύL�}
D�p�ś�;�*[9l�R�U<CV/=7�Š#��Q!�ϰ�GN�����P��@����_��ewv+vN���5�u�>���\�'
��A�V>��} KH�#뫪�F���m/��J H�Oo)ƛ��̖Uj!��q*�Rbl�Q�'�ɜ	t�1�G�I���\�`x���70Qo闩�Mۨ؎���=x�11���י��ؾ|M�Ԡ�{X�'xG����w�@�)5`P%2��5��/�޵�#���>�m(m 6��RDN{�DO�5�� �$^������A�<�.��s�R$�5�#Ti��1U(�H<S�7��C���t)VK�㊉)F>��*OW�Yl�F��B��v��֫߯(O����?���2N�F*��Ś�s8q�	8I�g�����8�9٥\�9����h�ӈϭ3�c٬83`�#�B����
�b�2}e%�e�8�,��H�hN�^��$��M��h��jv,|����4�0�,��r������?�_���X&�k)qh�3���?B7��<����pd5�d�V���I�-�&'��WC����jJ�)�O�B\-T�9�n
f��BA=�g)E%3���[s�/�-RG"+�F?`]���DVr�U�(24$K<ĝ�@��D@�<p�Y�� �F�D�`��6�ؐ��6�525]9����+�3T�v[?�aHX�d�������H�v|�J���p�b�Ytp�8z�^,S����OXz��Q�h�<�u8��x�l1��|Y��fY���;��,Ί�<�&�?~Hv�Տ�7I)e�V�K���>ȭ��h������D v�������S��N�yCU�J��j	�š��A��7i8��t��I�C�MjP#.ns�An��4��v%ԌnEȭ�*2�K�����R��3�`.h�r�۬��f��V�x���d24:�Z��]bUL����S���]��p~)���*`vkA �h}�� =��A��D�p_���9Q�l�#l��-9'�z��m���B��<���	A�n�QC��`�#���N�i� ��IbZ	�8o���G�}_��6^���c����Yp�r�x��8 ��+�����3���q�b�?xz�! \�V�'����t�:�H�����e�9�Y;ѵ?�q~�=8!�Q�~�<��D�"�FST]��>>5��Т"ox��E�Y��N�\�Z�A�u?n�M�I4d��%��Fo����I����!�h�e))�y3���Cyۚ4��t���tj�wj7-t�t�<�D�D���f�>y!��Ń�ԉr�����`q	|�����Ρ�RO�YGt��'r#Z�n�4U%�?��\�j���_�<�F��� �j���I	(˸�2��j�a(�yc*��6�m!j��M�?n�BBeD_+W����k���7P�C��'�NS��]�g��8HU'@�%,RR���͐|R3#q�,�縷6��+�v@ǽ[���k$3���iL��(�� UP������	�����N�?�`6�x�4�h�02�}����4�ЉIX�(�S�`�6Bq���fK��-V�w����x�ӷ����P���4P�����U���ј��P�
�o>n}^b�Ⱥ�̦Fph$"W;�m�}�9Y!4���r��~GQ��{�����G$Ce���-�a�nH�����,���[�M/���ڠ[-��&~��Ga�ڊ���oL���C��J�L���J�P{�L�v�S���L|���6]�B
�IiN��Azp)Ʌ�u������_- X��b��ێ���M��T:���.�I(���+D�|�����N��@�*�]Yv���"��E{��Y8�)J�Su_?+�����D�-�x]�һQn/x:��ZƢOB-���g�)``����a�؃�B�g#�J����It����z��J$,-���r�
�v��a�,xs�{U��`	p&r�'���_�Z xU�6<�́�����%�}%-��\�W�g��B�ҥ敼?/�.%ftnC֯����Q�3�M���ǒY����8.������#s���%�aO8�j1��� 2�q5�e��&�v��	{"�2��ߊ�u�?��z����\���_WE�8��>��b��� ����u�%�X�1�$���1�=�nJ:�|xT��+E+?��a`��D����&�����۸��UM˹!�	��{rIn?�\f�}
��i�]�B�����^:�LV���(�ϖ����Y�`
�=�d´2KDF��,�Pv�n�)��{���ꍜ���_.��� ;yж�h4��'f��;��-s�!Q"Ð��Eϊ_"��吨�4� a���#J��ې��Dp$�d
�lx�t'��x�����j���z�g �¦��Hn�1zDA�9�ɱ�w�3��!��њyk�s�,D"��U�!��"����Q���o?��A�B��H�L�L�LU��|%�O���T:�P�S��.���Ew�f0�UUx���ͤC~#iؗ���!�M�&��=��n����03Z�\�b��`+s��~W��|�����q�dĔ��D	���Ҹ��hp����
f|ژg��䆩�^��� ��0~_�ś�{���M�̐��e%3��C���������e�E(��h|:Ċ��x�A~�:״o3�G��Qc�GY�S��I%�P �LłO���Uϵ��,���F�u��cP�'�[@M�
�����/���g���6�+	�Q�eSȠ�?k	���9��V9��z�t>���c���`w�ܣ@f���j�x���U-~BhA.�ny�U/k��YG���2&fGnGѦh�����M�w�b�mXp�sC�)��N��O]K�_��yM���X+�)�w�m�r�q�k�߸����V[qd��괮)v�RΞ6��hN�f��?��G���p��#BTH���9�:�B�����b�Y;��p����U7ݠT�P�����&�>I��+����o�g+�ܯ���SW���k�D�[��QR�r? ,Az������鲵���ھ���v��UZ�!k ���C�1dԥ���ܥ�[��N��l�f~��IW˟�as����/@X.'S�!�6���2oЁ�n�IuL)C���f<��ӶI�T	y�ã�N���%���mˉ&��yP'��c7���8���L�VE�Q�q�1q�"/�e�ZJ��hQ���;7\���ֻ�^ȴt�80���YIu��;��h���#�sB�+��ʲ�P��s�M�!h��O���k@aj��x������Q��E��d|���-�a���r�R½�B�9����k��yr�u&ǡ���xb؃q��N<�[��zJ�٘�C�y�J7m��І���a6N'X��4L�kΓ��yjoŎ�`�1�R��UF��	W��Hd���g�&4Q�|l�v�l�!e��x�)./�?#1����]�5�l�[��v��E�lY.J����W@y|���K���������y������5�Ѭ�wb��sA�DZ�dΥ�լ+v�x�!Ȅ��e���K� �$j4�3�odj���t�Ci��I�zI���նYX
�ٚ?�8�z�)��7�.����4�7����$a����,k��0���Kɖ�Ί�YKZ�[]�'����a�H�'���������Ad�� �}�`$�����"��]�!s�T,>i0�UT�
/���8�m'QOd��&�ga]٤ ��_y��ȽP�i2�J�J	l���T��p�iM�ͨ��*���e
ag)z�Iڪ����<����~HF��ωp$t<��h�eV:�6�;q[c{��@�l�����0�"o��	��沆'���O���X�I��-�.����|P(�ʽ�~���-/��o�y����rKa�˴�?а�#��En���x��;��8��ʄJ]��N�X��-�K�D�\��4yV�!z"�F	9a��Fl*T)Y�����/h��M0�9%&l��"����:^�4M�?�%M�㙐���k��R7��2#Ա�=���C���N�Uetmh,�¼��M?�k�zׇ5u�M�l�6�*jB�ɕ[͢n�J�b����H<��٫%�ۆ�IЬ1o���CM�x�Vw�>��X�>��>k�������IH�g
�#y�l����~m�UJ����v�S�Bh�
�d�?�r���#�U.FmnJ}�,U���D�Q�	��j28r�c?I<nՓ,V�%'�Ͻ����F�$t��v��k� ���V��k��w�DxSW����4�]�� ��d>Z�nk�m^
�:G,������pU�U�q����̅^]ȼ���
 5����Y�{l�a��
a�:�'CL�/�^�S�81�\��R*�}��S�'��{d`�;�D��-s�M��j$~�р��L�� �&<Q���p	�D��$h7<i�lw�W��%ْ!b>��� a��Q]�*�:/�dY��CAy��>�h���>D�J���$�ڼ��8�r���'je��~�Wy^�|.h1�����3�vm/��c�e�9�ʽ�4�ᾯ�5�׿�H3 (���8l������n�����LI}�����ێx��\t1eL��+ۧ�0FÓ� �� �Y���Ss��V�����mpa�rSw��}�o�;7��O�.M����f �W���zN�(�h�����m��s�OB�'�JwP�y ����\w�����y�Igy0gʹ�1� A\�����{�J��0~�D�"�=��*��x`�T����u~>��SQ��d~�FY>��<2�Q龅l�Ƃ�v���E`�{�2�j���Mz09/=ə�#=`�32�L�P�@�+x���q3�]��qv��`-rD]�~�Pv�� �K�q����~����|���J�O����`���F~���T���+��{��u��D�Lw�����l�y��M�`���h�X"#��l�����0RsVS��
���u���a["���������� v��Q>)/Fwr�&�?�o!�{�$�j�3`�$�|OZD��r�#�>�F�M���f�g�4�9�0�Ѿ���h��N36nA�����a0��O0�N6�p=2)&O���=Y���9j��N����F�����|U䇽����爵7��p��G�u���c6$;�ӂ&�am��{�me Ӕ��T��/��p�&S1�2N�� �"����XJ��&>����qIA2�d[�i�Œ� Q�ͪ��;��`_�7���M@�+�׭�LY��vT-�� �hF�Z
:������-�8P�~������H�p�œ0��ܔ&$3USLR��Tqζ};��}��S�'�2�V4M�.�]|]�dɪ,MI�\�~?x)~Nu�������7�U^8�](�ّ��K��;+��R5���pA�����:j��4�I��f5�Y��]�|Q�V�L�����uCcF�Q05�d�ŋ�7��n�At��STP��Bлߢ��U��@_r"����f%9΃���&.7�� �V�/k�F�b|!�eN��_9��x}m�/q��)o��s�f>ê�v�9��ӷ�����$4�?�����\;�Q���L����}TZ����Ll��1֝Y�1_��0�y���O��Tl9MayN�Qc�i	x5�F�&�ig=uY.-x��Mt-<���m���!��`��Z�A�����;`$^�ݨچ�e�9E)t���Q��)���aZU�b��1�mA��$�R���*w�D��X�5�ӣ2К�cϠ�T��tf�K�r��OQfwd�mgƷ���1��k�2f��i��l��8��� Gbj�aKZ�5��d➱��}x%I(�&R��I���-���I�[���������x'<אAJGK=2Z��זG�̝�&��x�P(���sҊ��ͮ�S�E�ӑ:�%��U�b	_u��P�Y�WV��8��a�����H�FO�v�1�@+_3g����`'!�����A�����$�e��t�aW�;�n�4c��&�㴡V#�3��z�m�AcW�Q&��AP����
��)9t�e�������`@�8�Y���}��R􈩂�s�� �N���N�o�~���.,�{����.��&dV�����"�	�xU�4t��;��`ٍ�?�:N�Q�u���ԓF@��U�"]�KH�̹��s������ ���b��72�pi�w�};1F��C������Rg�4op��4���X�G-�
3%����� z#*��Xl]�wr���?`�5)�u�_E̬FB��w����i����$�h:Q�6���<�?�����`/��g��O,6�� M-b���V*����^����/�NY(yLC�%�ul-/0mU�b`#(�f�a��J;����鄛s_�*4��\_�j: e0&0�����os�T�j���B5���U��~�m8�d@�����{`v5��w	�|Lݟ9�|�=�C+9
7!��| ���&�>Ih2�臸�`?{�g��q	-�=c@���8q����F3�0@�x�d~�¼KQ�}8]�=����釩@�Q6ҩ��R���;��s׶��r�˥C��G��A{&*�rAe��sp'Y����QF�.ػl�y48.)�������T���������H�a��,�j��NQ;-�eRJ-��-��c�^�Q:�Ti��g��_�c<P>�tA&�05����Yz���ay����5*��\0j+`a['H��&ԬZV���pq��i�t��şN��s��$G_�U��ys(N7D��u<%�X�',К
�8!�	���Ű�DP)'� s�s�p%P�l16�)��Eڼ-����G��lS�0Z1����:9�`"C2E'w/�^��A���JO7������^��������p�U��?,���OZB@����<����^��(kRgw�}&��i�H��ZH�uP��:n9Ϩ��J�בcRuJs��(ա;^�@ �Ш�Ę?���&�ǝ�$S?Fc6 �+6k�{
���|��j�X�T�M;U��lI�T�i���׈�hC�y�B`X2�h<'�cpL�W�'RZ�XtK�g�J#�`�!$���#GC�Gc�#�✤��m�	���4��$��u�/��"xB�}ntc�pH�m3�)kz��4n_Wa9�=E�	�}��h%��TT�R�OҊn\S&����:W��ᴾ���X�w���s5ݐ����WZ)�?��YO��ᡔ ����]��N�~�CI.��4����K!�l�l4n&��'1�˵�}� �,(�C�o�xQ~zZG.L}����ޱh']G��c��|����G����}s�>�$���8�%Nb������4��/�E4�AJ.8�����7�P��� 	ѝ�X/Q3c�GA�ڎ�v�2<K�V�sE�����ļk<� b�J�Y2�"�����<��񡡈|� �%�U؆n�K��L�P�~F�/�Q�;Eq�d����=@��W�R\`�N��!1r�*�t�<3�{�EeC�&Ԡ��	�Z�Y� �-.R�_�=�����.ƪE��&z����X����*�G��ܢR��"��S��i�W�!a��ύ<q����,q��7���Ȧ�̲�C�����I�Ǌ� �<h�C2��1��t㯫v >D�􆝔�z�3}�a�]�R��O��}K���6�ؚ����I �o�I���oT[�͖߿�Y�	wT��<Kwe��ÉU�z�ޕa������*F��8{���-�^����Gx��&,KM ΰUVfhvO���Y�}ď�������xzc�:�m��W*�_%�܌QfPyym��e��"~�猢v�{Ci����O^rj4D����>|` �wv���j������J&��8�~�����TK���]�F�L����߫v�<_�w�Ư8l����Z�����/m�^�����;�r�����2�P݊$o�Ȃ�{�J��!�J�i��'s�t�%p��Y��y$,+a�p�0�#����z����
C����"��A����9yi����m�;z�֝�h8�{������M��Q6�b.�/��*-O_N	p嫩�.-J��e�+�Aa�h���V\�xשׂ��Z%㶆A�Tr�d��4˫V��Ѩ�~$G�.ku���-  ��c2X!��r!�%�4�n�ǜۡ��!"}�XꐒI��S�F��!�q�	_T���,��W:��� ������_�@>�k2B�܁q�+/���sv�&}�uD<^�:`F��[�-�o�m��gY�e|�����~��8�zpk怢��7���J充\�r��<�^r��¯���� �>����u!_����~�w�a�ݣ����\>���u;�}�MR��j}��7��讓(�^˿�ǽ�D3�V����\�㐡1�J��9���A��I��z��!�^aY��:4����拏��
I=�7�RN�{"���y�jV擁�����	H/o�$��:�`��6�eU%�_� K��ڹfF�\�5)��g�G��@I���?:r��������/������K]G��W~�e�1�C��S����39�T�?O � ���(�l�s���}�X~|a��3�,b��o��	��=Gcq��\k��#�}�y`��׀���B-�Y��B1�DL`�z�x��`�%r����=�F�j��P���&���jY�u�#eΣ1�70~���8{΋���s�Y�S�1��=Ӊ�M�h��7<,}4��v�'��p���tD�&�V*cm�NVF��t�À��'\ �;��_�ws�=������D�w��u9��O�i�_��h)hq����|��l#١��:w����\���\�j�?��tM铌��� H�s#}�dM+CΙl�S�����/��' �(Hu�z��N��e�cSlߞr������`] -�Zn��6S��]����Ao�����{��]���Z�ᣮ�Ṽ����ؠ�x�l>Y�s翿U��<�z�)NzΟ�=,N 3{?���ϥ8j��Gw�����[����ҷ�9R��n����X4��'�>%����9�T�#�v��9=���zsx��wK�x8����N����?�Ӎ\0u*�z�N�%��-r/�۩QY�j�V:�Z��p���j`W�� X~ �xa\K�9'��b��P�u-�v�(�����p�>�J���Ş6�EK�k��9�6�*LD�N[D:Ή�;7��)y��VP�5���)ܘ%��Hl���	�c,!��ʸs�J�e��q���vZNR�}�8H{T�ƹJf
Ѹ)J+��3Ae��3��P��u������Qw��$j	aHD�i�@���SS��|3m��vY��iTڀ�Gn_�;d���S�7.E��_�%]�!pg0��Bkh�W2�Ya̽���F�'3���	]Z�k�YZ;_�˟�F@+��j�ʁ<�S;�8����Y�8��]qY)Q(Z�W�poO���ǐvW�yl�@�����7 ~��<�Xw�$$����\�4�,��Y[U#�_�P$`)�ǅ�+��`����
�T^��9R!�(_#؍��G��
����j�����j�6����^]�̐���U8�R>��-�#�3�8�Gz���Or��AY����[������e1 ;�(���*�{?%����M�g`r�G��Hg1��=� o�z:�7^L�ϑ�}A���AMB��N�xr�`r��\�:�iаd&�|G�|=�'xb��n%V�&�Fkpl�El�I�H�'��͒�?��8��.�kV?I�U@$�P�v�����������!B�8�믝��re{g0���`w#�6[+�a8m�=`�շ٠=��f�`��*�"KL5�Ͳ��p̼��}���.�ћ�
B�-��Zu3��tA���:Etة.�1<�� G��r��R�@-۬���J��>��3����?�iY\�C��F��o՜��/�jC'�����ʶm#S8y!]�h�}ajͭ�ڨ�R�2��������X�;�vp��9�����1��ڈ�����R��������M�8�6�ps���W���D���k�p|`)D����1�k�6%�eߠ�f����&1�g)�(n��� OtH�w�&Ux��VIQ�ܩq��� v��aUk+��:V
���w���,�;�̦k�Ĝ���O������'U�� -�p��bD��c�Th��IJ�x�&X�;�PzDZ�\|Mt��m�^{Z�'��|��0[�Y�ۻ�ȟ�ɚ��}��D�&KG�ѯ��Ǐ��,@S]��~.���ܮ8"ev�!�ݱu ���{�b����g��3���g��/4�� ���Uq�N�p)�{t�]�N��E�&A�t5 ���OB���/=ck�H�m�ȧ�&���e EP�|��-��zmK��#j���<����f�cVn�_��;��O�%�pŞSD]��X�;���T)1'�T��n!��7y N��̼?�ɇ���q�����y=$�l,^ژ���(/�j�u�rҭl�$�	񌰀�'S���n3���+z ��;����xS瑶m�u���^!��l�Bj&&ݚ�O��m1���w7�]��Vz.ާjL���� �r+��Ӎ�VK ��7�}�16ZY�Ԗ��� �9�q�
O��4^w ���i����Γ��_���(������}{� cz#�Z�'k�����zϽ����9<�g�������*P�5V�W�>���=��w+�f�n�Ϫ��(� t_�,��W�����5O8x:����arK�i��B�z�ݨ�*Q4m�+]��B%2՘�f��f���o��`��t���g�4a��>�����k	�t�D��0��Ɖ�0ތZ�Mt�͓uq�csk�u��Un���"I6�!�e��������i%�I�M��a�:����+K�Bb�Tʅ;�?j+YĆ��~+I�_�!E`N��I�3wi�&_;� �tfR�v��e�����ś�P��D�N}�ѯ�͚��Y�Gn1�����'��R!*������2~Jy���$i��}5��oPfU���i/yքp����Z�Tg�"U�O�o<�d��Xb�ʭ.��6Sk~��F��l'�e�b�Vuו0��_h��T�������:R�d�i�ذ���݀��r|�4=�47��3���������-��5�s���,x���� ��D����e�(�^ oT�- �����T0��Z�?I��T���Nj�q�ӯU�0r"�z"���A�B�;�V��'�Y�w>�����x��	���Ԝ}ٱ@�Pj=QI���ob��Jw��v��9b���h-����:��V-�BE��K��:!X�
�&�a�Eü�埶<sY�!� k�XG��'���T�?�t�Ӷ# ���W��x�?`:���.5�w.`�|�@ضM����!�jEl�N��s��{t���B�V��~l�h_�N�k����)�ŉ.�f���z�Ѱ�?�X�ׁ�`m�����Kl�eX��7�A�*�SSd jc��yc���f?I1�mI���m�/t��7%Zvf�n{�e#�E2V:g�3�ǰP���7����[�&��ց��p�����x��s����[#���O�,}����z�R�謓$u���(��~g���+�����$��G^PHX�� f%�r�����	b��.<�(A&t�f&9I
	U�X�'J_�m&T}�,�G�r���,K����Ǒ�5�(޴�l��D4�P�����Q{6t-��a�	�V����^ ����0G[�i"�HG��c���K¤�x�~O�e!K�^ܚ>)���&1��7e$�i�5��)��M!��w��Ɗ�[3kR����Bu]��el1ߠii���9f,x���8�r&��6L$��GJ�ާV+����c&��0�7��8��BQ=Nf��5;�8��qx���?V��rd���m^��+�sE�+ۉ{ǲd;PjwOB|����偂��ZXn
���B�6�-�F�DG�(g�/�����p��sVOS-.f��evG2)�"�.�1u��Շ� P����j�C���V��"A��5�w��Eyf,֙��K~Jy~�o(��N��}��u�#�4 E�L��;�����G���,��Q�Xa���|v������f/�CA��
�:��rA��֌�ax��[������\瑆��&�*����7��B�Q��M��\���QqÚ�%�"�F����?x��G
���>n�~6Q�OH�Y�-�����K���Hz=<z�D�01-Zʔ	�@Yx���i���dy���������̧�ލ����7��U<g{@�v[�\�!RpCs#���f�N��ql�Z;���Y�|}�Lڊ�Ń.�q���/E�|�\���5��}�g�w�!�)X�xa�+�B؉�4���97��6�#��}�!H�xg����P{���t������lnSka��t����B��ƈ7R��֡��.�d,ڡ�(�F���T�r"u�+z=b\�V��0�/yK��k��]C�L%E�
O��9�]�q
���dj�)�[�JЌ��fím�M�N"G�'"�,�Q\�l�o��Q�/bEJ�<��鍆�������Awz�vD�by3�V.D�(�ZW,0��C�쭐��������9<L:�h����9�2��c�ʤ�۴��L��W�����4N������	�a��#��$�3Raw%з��gj7����� �E�=M��
���&>�i��"y��dnCy\}!��p�m�����b`� ����~�}�[���z7
~	�H��;�T��Ko(a���!m�E"�WD�ް����;����p|"-]K�?Pv�rI��)}�q�N��X�0)�	���zk�u�:h
Ŭ#d�BC�S�-06E/W��t���(�mMP�)U��ե ̤w��L���|�D]殞�r�n7s~-�g��i �}�h5���y�~�9�����p�vm�w�G����|�nAp�$w�~����O�NZ�,X�m]p�� �w�}`���큛�Gϕ� jP��U��^�o�}�/l97O5����l���Q1B�Ǒ�ސ�W˵�u6P��j�Xt/��(�B�g�C��3͉�%��g����;/�l�<=9�R��Ry�>����k@E�3�O9��'�%��L�Qmze>d�m,��W+.�Tm{�5����lƯ�+\`P�zhju/m��bc9*_�bQ�{ '7�pOe���c��9�h-:�}A�b`	����}�
郬a��	�^�E�t�hJ�~z�s�:%|7��l-�*���zغ�.k�!#:a�H��}���u,���ۯ��>C�cH�:��q<���{4�<��_�qkf��|Z���ow��@w_Jx`��ڤ�y�̈$�L���[4��1�Y�������� ��E�~�	�ط��k[�+��M~t��0��8�=O&k�[��\�	�7�OHSI�=G�Dd��	���0�~nS&��4�IX��4�O�f
��������������(\�K�Dל�8��
�½c��i�
 "�>y��]�������i�u?�U_�3��-��sM���'�.T�<�"����V�w��T�1�c�H�I�js��dS�Mam�nJB�K�(�}�6��/fbl����Va�\=�k�E
uI�J�A��kB���'�.JIrx� X��$��<�|�m'��rr��i����X�Cv�䏯y�$��*E҃��x�<1�1Y���x��-�a���V]Mw�J
�(����7t��$cr`��0�@
��7����z����<sY��
��2y�030r�$/��0���镤g%NmO��l���@��Pj��B{,�_rN)l|�S9'bs�$oq�������.��čab�Q�Mn�&G`]w���9�v�~OpM�o��ٽ�t�d���N�T�p��jH$y���<?���l�$�����u��
̂Sk���a��3��&�K刷Î������_�[�+c�%�W�_�	�+)+�>z2u[AEEA�_B���NI�n�vn���g�n*F�8��ƈX��J^O"���|��|I�/�7ÿ5�؎���{� j���zt�)�mtm$	�N�A��y|�����F�_���FfV�m�V0���LQ�>h�`{�Fl��Q��%��߯o���l��(�&�［��6���h��3�A
�~�������q3����&R�<��Q<�1�@���n�j�F� �JM�x��s�L(�e��H���(+0��QD�j��7� �X C}y�֙�4�w1�\����t�۳�x�y;j�O�1�藶Z@"�ʴ4yo|�r�bl�>ԫd�j.���_{�O]���^���zdޯ��,D���*wB��5�wh���q0�	�ɇ�U<Er�g�jX��eK
e�k�ݾ8?wY�ЗE���1^'��A'��- �iqtȦ���4�C}��HK��Ef�W��YN$��|��f�1���9���3l'>�9�J������k�+q�!`/�J?�*@����T���1c ��7�6�G���gI�~�.IE���V'�Pr7��-1m�!N�¢���_����f~c��mk0�!x@L]���'jU.��'����/�`/��_��'�/܄<9L׸b��m?Z���(/X�צ���'C+�R��+TR{��0���~�eڀ�+ML�m�y!«-��esZ���&���ȯ	ݕ�_�\�8��[�Ec�uC���.�b�oS�!l��D����TD����&��Be����ʑ��D�T}a���`�U-�9���Pq?���h�}�l�ĸӭӨ^�W��I����5�|oZ�ԁ�ϔ����vO"^2kY� �k�����A�b?���r>�-���/2�D�- ��Xkź:�Qq� dAB��,���Hɮ����'�"@R���q������_�Y���������FX��"�����[G"q�o��5\��Z��dP�p/��K����qc��z���I��ಡ`�e���b���W���5:bÇ�}��=E���r.wb׊
�{���:�@ux$<[f����~� ��ND*؏A�.�b��#�ȡ��w5{%=���+QA踆�L���_��1���bx2�o?iL<�~T���cpp��E�^���&�zi�p�9k�ɘ��
��)�@�`����Na�Uc h�EG�h ���0S� �<y��2����y[�Vw��KSp@D��)�}"~��z��tn�IjE��m
]�[}����C���e�g�| �!�fr<���s�DE8j�V�DF`*�wg�D�|�D�����f/��f��7*�=*Q�~*_7�{2��b�#���'~�<�qx��ŀ^ӟm��s���m�_\}y�Y��:�O�N!h�-�v�d�Mr������\�\{U#@D�d�LJ1��p�BxK,�|�������i"j�BH���"�;M\���sl��|!�u���lm�O�qś4�8�X������H��݈U�����RG�ޣ8�R�eOd���
���Dq�ᢁr	�"���~�/43?����~��W&�4�F���d 1��<;��>�}�k�-����g�m�IQ����Qa0�p���(|�	6�E������d����G��)4�-�� ��<���*Vj���A�x�18��Q>g�)�������3� �pYnx���QK��A<w%�כK�A����:�^�_��K�ՋN�t;�{��̩�aY��iE�Ii-���}��i��]��P�׵G�7/�1b�^F����%��U����^b���o�:<h�=t@��6����	ҟ��b3*�Q�!;��Լ[Ifq�勅P�~K��w0�<��`��|��e���e|�p�c�B%��`���00��m��W�&����q�/��(;���5���6�)�����F6b�h!�b����@)T��)-�:�,�ͥ*��JS�S9Z�?�����&ug�ZV�f�k^�5.\v���Ư�T�r�#[���i䄗��,���2� =��[��p��v˹lx��I�j�xea��CJw��c�� δz���7��o=�Ȼ��H��B�t�>fN*u��$�y��n���{O/�ݛ��z���F'X���Pj��
$|��FJP���:�:0+��/ C��lφ��R:ԕ!m.�w����@�T�jI���^������9�ihY=�v�����h��lJj�r��苰}�[Q��Axj5J�o�q�ԩK����!eD�2�>�I����W? �Y$�}S�>�����8�g<��}��
�D+Z��͊M Q � �7�|:�1]��E[�� 	X��x��8���/���v�iM��I��e!b��qb	�C��aɳ� M�8�1���\Y��Z�(�%��A/A��*��>`�b*| �%����D��g$<�8�{J���Ft�Fy���t\�(١��1��=؅.,�p�ڬE.����cT��*;�F2��j�A5@-��Dr�@X�0q|o�"�9��u�Y�vl��"-��?j_%/�]|R;m}�� �a	�bTr�Ӧ%�?&þM<�tx�N��'��Iu���f�̼�m|�B|/T��
%(K0����;?���g��{h'�F���3�iȰ�����Ev��LJ�E���!�?0�!���92�EO�~���K�V�ܢ��~�[���Q��\o��uf=	:�?�I�����v]��W5��o$	��[8�'�t=q��Z�I�c�	%���i*y�4W��*�D��^���S���j͖!m������rě����ȓ܋	�
ĩ����ir�C.�.U&�1D�x��)�������Y�y�ˢ����١�~�׏�'�.B=��'���ӷބ��n�����+�������s�S�w�B�����xL�:^)����ۛ�-�ng�����s:H{GĶ4���Y������C�̞���j�K�9[�U�o������=0_.�V����> ;'K�ar�T�D\��2����d��6cQr��d�U�)�HQf���>T��Ev�GS�MN0����Pb=�jZL�"���s�
�R�_:���I�#g�����#3�U7'�V�����K^*�[�Iq[��
f�N-!�)�$M�Fb:�]�͋r�^�Vz�jb�ՇRD�t�vFE����(�k�By��E�� L-�a?`H�!RΈ����3��3���)b8��Tv^\+�r��^�>O�䃶"�J�;�T��]̮8T ��(�vM�����WT�D���R�v�
�4�z`.Y�g3m����O�nY
�A��"�r���(�.<~߾.�-ـ���
��˛53U�W� K�Qu9[h�B�����kv�j��pf�קu����W��h�/ah��P\��״}���Jf	�4nLL��1��#�����-<ni��ǚe�1��ʼ�Y:/H�8Dz�T^Mc��	���[]|(6�</�0BYK��䝅�����0m���u�<E�9ox��r�54�f���gIO�|_�@�Ng N������&��9�-��K�nԸC�E��+o�4rV��C ��TvS<ST[��N�u����y��7���;��s�<U���A����x�,��a���@�!u#����jbE�Ԡ�a?��Ŕ(��C��u��5:�&���sG��1�	- �[���R�҄���^���'B]l��@��?���V7�/
��[%Et�{{�!9�L����b@Pq����j� 5�4$�zKK��H�a��CV��Fx�l3A��B�G�N��%��RL�Œ+o���g/f>�V9ڒ���X�F�m"����g�	��{ĢD�>�4�/�"&v���yh��� I��;F�D���,a��.�$5�5�)_#*��$+�����p�Jq��m������
1�Ȁ�y���Nq�-j�S�����o˪�:)��$'�cR�LH����{�'	���Z�l0
��o�Rbj/VSFL����C�j~iSJ?��QەI�7kg#���+QR{X����|v� ,A�C8<V�g��8$�]�E����ǩ7�\���ą˒he_��|ώ��q��i�|pa�8XS�֦�˫�	� <-�nȏ��y��%?�PDЛ���q�^�?��1�d�@!K�	j�����Rt����9�E��YBFBK����`-�}a'��bĳP�چ)δ���%��u��w���H��Z{���� �v3��5A�������~v���Њ��VRM��g�j�1�z�!��"7T�a��n�)TE"m�5�fv���^b�׵��Lo.��~�V�N&��	�]G�͒��l��[y���es�b�6P��X8=3��5��pn#D�A1����#b��)���s޹[�\ �;PPe��P��A�ް0N������q
=�������͋�gɬA_'�/!�Y�YK�!@d���!D����p�����@����Y�)���B ?��^D�iՔ����4�%�\>��sI�
����c$��a��?@�f��2���1�u^���=܎�VP�"6��7�;֖�ZZ9��ۅ;���i�ȖKɸ�ƕ�^���*�ڄ���+��ҶKW����s�n��$d��}��z��o)sv����[5{��z�q&�V-��-��ϔ�D�7P�e��V���lM(�!��7v�%DWY���̮y`��I[P��ɱ����G m��Z<%�,C�H���^��7<�P7��������d4����m��M�AL����Y���`��m���3t!2(���Y�d2�������_�������	,5u]���F+�z���M�:2w��e5�x���7���;��|p�}v�~���p�	���qY\l)V�,��&�y����g��<G���3�B���P�� %�U,���^���b#Mߠ���_b Nz*E�m蛕���0�䘼���v�?GaʽbȾ<���
�ﯬ�x�qf�Z��Ar�K��a�~}�m1[��]:hZ��8A��U���V2$��)�:�H�P�3G �8�C|蚘�X�9�]J�|}@�gPJ��`|{'J~��_�vs�k����^V�^��Hm���y�����S�\ΰ�6-��/��l�Gw�فvCpH.eP���h<���H��w�Gǩ0�
OM�3ißyt�2�eݪyWZ�r��t!�z�{I�:n�u��l�uL��[���(i}Q4W}4���c)�洞Y.`��am'��1� H>@�~�hW�=�L�E�����C�?`������r�/K�ȗ���ʚ�%{�i�7_�qk�EUk#��P@��_�)X����v��R`y#�f�7$᫈�֌[j?�������S�!�m��?ܑ㪔�}' g�Y��Xy�F�C���㺈��57#i0'���=���)� �$��k�也���N��㧙Cd{�F�֐�~L�u.���t� \q=�6l�@4v�����`6K�7v`��*��׼���^�ѝ���,ǚWMqx�T�?7RK�ys���N#��4k�T���u+�����kO�PA��y����Z�P�)>��Q�����\`t�,-"Sz���=F����50�S�[H��%�@s̳������aC�Z�ޫs��W��2M����r�y�e��QQ����y�a������Z�Ɓ�I��4�'jA���M���O�bf�
�]�2ɛD�6�o�J�:�Ra~A1�����(�eY4�'P7Vs�!q��
�"w3�Q�����_��#�����01>���o �2E8F�	]-),�3��nx��3.��� fkR��,��N�dI�U MF��0�����-�,#��,�ɓzZi�@�6�-�1��V4��Z�X��QxV������{\+7g����%+Q��FFD���Rn_!>f�p��sPB�"w�Z������W�q�X��6�g�˸��ϾHh�wTc��L����i��0�;��Y�Ø|���A,��e@�:��f�=PiA揞P��8@	�0_˻u�R���5F��5�(f����*X�I,���+��I��p�1��Uw��?G��������Nm��OQJ��Ȫj��<�
] k*�L������� �J��c�hɃ����^B�|���%�#`SJN��L���a�m�¯�b6�Q�ρ��|���z������Ω֠#��?�Z�1('rBn(���̹�U���$�h� ���'n(݊�t,3�҈���4G�5�gP��J��򳩛}Z!��;O��k._��[l.�[ڀ!. @�c8zNܕ�n�,�%��Q7$��R
�y&K��O�e�����<�զ��� ^�
���}����f��"���n���Q��?f� ������%$V:����pV�I��I��:ڎ���Va�1P%%��g���x�q�_��A����K���_\.���[���Y#'4�L�C^DO����Ȫq�>�li�e��f�^K� �a�=A,�_�;t���o�>o��C�����?��Y���y �VG���Q�)�Y5*����7�	�g���b�)��
(��]Y�����U�*�lT����|N�ܯ�H����d8�ʶ�~&�*
���,�mXJr
����=tA�2��o��,z:�~�X�`]��|!GSA^�a���`�@v��Y|֓Jz��_��Oz8�H�ǔ�C�y�QD�s�FN��~����$�0! IB�h�Aj��d�G����7U�� +;5<��!��Z�{���s��"ݏ�}��°�zA�5.�ۺxds��x�ue�mN��N�E�6nxw���9��:�T�Z��/upٸ�Q4Aڥcl�E�>/�)�J��+� C�!��j���AsHy�ZG�}8+��?|`n����Xs�����b��2s�
��j��"���=��!������2�'�O���X_�*�VQ�ɉb�S(%�l.O	��(�b�jV��?�� tM�@O�C�~�*��%9�Ť��վ�U4��� �Q��'eN���!��E0�wA�Ӡ�E�U!��)����m���	��>vnT������A�a>o�D>�!���l{�j���=�8Wb3 ���}Pp��#�%�%2HN��`���U�{�s�������b��4��7�SoY�p��	k��e vn;��3�P6<�Z�X���0�+{���ّ$�t��>���3Z��7�$�/���Y�D�e:�:(��R�	�W��з�ѡ��v�v,�Y-9��}]�6@���&��>�>
�V_P�8�?^w��/�&96�ń!-�ʎWy��s�}a5��n��BU�F�j,�<p���d��矷?�4�{�L_���1D,`��t��5���_6}���BT*�2~M� �YMa��Lqifޓ�b��F���L�9ʂ�oS]�A'k�؊J��\�{�&ۺM$��|��UX�����r�� �~���s6K�+�����Y3˭늓U��y!րQ�60�y(�/���{�%I[h�*�+��cs��-/�>@*:��__��e>.��T����!td*�h(���<C@ cdP`Vz#�!�0����o�JH��0��`��������"C؁>^	Iy��T*����5��#�ݢ+�����?��IRY�Y��*��]�%u�0�^~)ʌ�Ji �@���O2�r4�A�!�zp��ws��a��`av
�0��9dh����_
d�70[!�b��F��U�ww'�2y�~3&�S���q�:
��*��7I�(@"���D�����)S�;�R�qԏ\Y2�WM��w�\$���v�2G�a��ؼ���b(�NF��a���w�3Km�ecG'��������F>TB�X�2��Lkn�VGf��бM�� R9L���R���t/��h=�D�I
~n�07���+n�a��3֗[��{�0�Ͽ���r��m��Ҳo��e�m.��cS�M6P`s��NԆe�o�����H����/�w�aD�`���ي�:�5�X��
�B07
��='6��s�3����9���:�+����~L=� �fzc'���vr7hn���[i}���j� n�)�rz�2.�	N�f2�;шf�	��O#p�o2�ۮ>�5�v��Q����8&���De�P3/6 ��HQ�Ԭ-��#*`�]L���QV?O͑-��4�(f��N_�7�n�O�\��s-�[�귿s'�j�lb͜r��v���U�F�e�u��6�y�i�s�W�~X*���/:u�H��4�����)���Eu͉q�ɡ%1��בCB����
*B#�zX����!ս6�a�P��Ft���=����AL��ӄ`x4t;/LEt�9��cO��4�C�{*��I��a��]7>/�~�:>6nЊ ��
�&<l���E�@��Һ~�Y�-g�Y i��r��UA�{#B1���x�M�ɫnO��A_.<��X���О`������~�q4Ɇ�Ɂ3|�%�j��@\�h���9��{������f~�	<�\�ʑD��h&,��w-�!6��(��T�O��S�N`?:�W��M�����~��h>���Po�IOy��Ҵ6 ���e��x�|0��{�N�±�&�����3p���?^M���&a������8��v�� ����x��>W���7�JN�b�%�r�mʀ3�b
��7o�ǘ1�ȸG�"�@h?g��X=YY`@�i�!6��7"H�xF� ��Q�ZV���:��b�{>D$+��dP���	[�l�k���z�����%Y���{9]�+��'п��ԡ%U�b;�<v�"M�_�
����1�(	&�j�d�����L�b������6ͪ��*<m���3`��{�F���]�8�̣%gTX	��&��y����C�E+����0/�ą��|��8�^��{�rO��!��{t�$Ƌ�v繭����RP^m�hD�����yzK�1V5)���2)�� w�Q���*(Ę�-�$�1��ζ�M��h}g?�w�_�Kp��|H����W�k3��S�6��O%��iJ��H�+�$���n�Q�!�h+Ǻbs��Z��q��9mR>ؽ�,p�Zj�Q��E�ku�����l
'�'"�$߳9E�p,h���OA��9�!�-n�z���A�|���»�v҇���pM��z�L:ݻ�8�Y�'U�V�c�#>��G�Q�"Y�����;����ѧ��0��.�_1���qLo^�ex�����űQ�9��n���(�ו��<��)��,햫�ڇZjAa�0����F����C�]��%��i�!%�gҹ��xRB��g�&��f&䳰��C�(W��*�4��SL,��	*Y��{bޢE6��вcj�Ԣ_; )	�I��L��2��w��/�KS�|�es�3�Z�ia1,�6���R]mU�)�� ��D����g�2�8f}�@F��H'$��|���q��B�0c�|���#���x'����Z�q��>��)�c[�]���Fhc{ʸ4/<��kƏ�rԶ�~bD��ձ��(�Π��eʤ�b1�~�QK�P+s��p>�t��q@;�	0FB+�p��"�@�����W����p�B��J �U�)�*����3���y�["XVDW/`�:7ȍ(7
]�k�^�	o��o��Q��l��.wGKh��/p��$!c{��(�b�Cb!�c���S�� �ݚs7�����C����xl~���F�d�k�3��h- ��p��a4T�K��RACURD��d�-���L�{i�cHimw���<Ce��G��_�34-�`�6X����S_�2Fƪ<�<K20,�Uk.&�BG8��_����޶^wwI���kҴ��2������jeM�}{�.������%X��ȓ�d�͹���l�s%,O.~-�5|1I\��vE�,nl�rm/Ϛ0�#�9�J�j��A��X%4��3?:����Ȼ����Y���eR#}Ծ�՚(�B Ŕ*��%#)���~�t��uL�F�N]
��@�@���۰��h��@Y��ؽ^�Z�m��~�z��l&'����4��H�&��Jx�e���P�'x,H�4��?2���[����)�8�� �fg�[�W��b6Ɠa]|�+\��
g��wW%���l�ƞ�޳9~��+���w�B]���k��G�g{-��*�\CH��"x'�C�<�����j��B�C}'X�D3��-��EAq���^�歰�bP�Ri�$��QɌ�T��U)J/���f�G�ތ&�J�.��8"���i�Gc�S�x�*�	?��z������t
�'�<G?l0��}��DcH�nK�7� 5�W�<6ה��aΦ�g�}��e�U�*�A�?�P��w����n�NT��Z���n�L����Bp>�A�sV�*4��w�S��.GZ]�:`0y8IJ)~8-��-�2�#���({;�93q��0�R1�FB������|�ņ[���,u�L'���3�{�S�.�`��h5T���Ee�tE;������~��@���P���M�{�)U�����,�!z�x��FS��g��(u��~��EmY�ա��pM�(���<7�3�@��%�#J�|�=��6.a�\�[$P��Y��ލ�����ˊ|v���UW³� &+(}�R���X �^e�]��sB�\!Yr�p5G�+/�5���K|��S�W8�9B�v׌� �3+Py�jy+M�M^��E�1C)�:.�ݠ�^	جAƈ�_��Ѯ��A�� ��j�hZ�%�/z�R�ߚ_�t"a���>�mC�����Acv�A�y'Sc7բ}6V{�|��TY	��1�/�vL:�S;tW�~�=MľQ_�.�\�^L�y��s�����܃	���lz�2�����`�}������F7f�h�X����d���U���G\w�˨��`��r5D	 fU�ъk*GL���X�l�{�ns��ز<��%�_�x� ��-�4��Ju��2���g�G�mr���Ђ9z��)�k��tr�0�����c�:��){�5>b}�ռ��� ����Hl�v�u������e���J�#?-Z��q��f]�:P���Nr6�� \Ku(��'x1�uFF`��1�%!�e��nA��`Xy���ٰ�$ݴ���l9��������\#6E���f�}%kr���S��������#�DnpL�M�	��`�d�A	�i���5�L�t� '�M��,-�E��첯Ǌ��B���6v� �fO�A ��@<�L��Ox�D����i�Ph,IlUtG��5��/.�(;SnI�?�e��r77{�X�^G�5a$�9�Y@�/>���~e\\)D ���^�x��w����kx����#Z;��jLnc��s8�­�H������I~��$�?Q��S2��,�`��0�X_�s�հ#D�[�i!$55�^~;Ұ ?4C��wx13E���ݧ����
�)ݚ��p���e"�
�2����#B�FՂ4�����A�N��f�����y~儐�i�RW�w1�O���m����:�q�%:�N*eY�w��]+�qlJ��%c���������e�!^������]������R_%�I!L�x��@a	�fl�{v���G�n�2��=�4@{:�b�@�ߖ�^8J�hT0��'ZMIcH`Y��	�T1��6�G��K?�v��3�n4���^8,�3q�N�9t�u�<���_�#S�K�m���1���*�~55���w������u쉏�4R�:���@�P���S#9��ƯÔ��=;M��,�!�˰�v�"��e�s���S&���&���#G�S�Y� H������iS��5��{�w�\E$|�H1p��ҠF;t�Cc{�ZV)�H�7m3�_�{�6�>�-�z�X��q��-Xz%�'�mK]���s�u��x�:���Y�٪�����Bq�_�����=G��C:�F�k�)ÍY��g�}Jm���_q��0
̲�k���k�p���/�"x`��W��Ώ�/i�,a���cK_��x,IO�i��B� d�)��m������KF���7-+4x�
:�ף��hX%E��% [��J�0MUOS����2<,�Jef�3-�-k�(����v��,D��- ��S0�C%�h"����3��a2����Խ��a�8��]�p��l�	
8�6�&y����fT�h61b��|?����d�OI{�x�G!�F�e۬0�k�]���0#S0k���_��甃��LcV�M��O��+/��U]���E�_ �~���&Z2Նܶ���H�=��!�C�Lzee�D�tRȲa6�_g͇��-%@H
i�ޱ��LR�t�9�o�%S�G�U 8��g�� ��_��Q:"�qf����3Ѐ ��I�kz�>�#��XK.��[u�7�&,g. C���J %��!�o_�'`l���y��>����D<s`_4����:*=fY�*���P���Um6���gE�2�6sy��|V'�]c�k� ~*�����}��Q̟q��Ɨ!�f��A�������X�[�g�.j�N��)V�cj�ɻ�;?���˳�l�-T7c�ݼ�E��^�����g�VOn�n�oĔ�������wP��g�On>љ�z�|�3�$��2uxCF��� �����z�W#����pϏ׸�?�����c��='	Lse�}�R�m��-�YO|�j}���㨋\}��v�}�����ݧ(���'�n>c	�[#�<�Ǉ�$(�#ġ���w>l{��˵��IE+�E�,K�nD �ՙO{h��D����~?��[W��4���踾*~�"Pˁ�[+<�*04�Cq��vd��K[��5�����},u1�B��YgH�[���P��ȮpT�ح��oS��~Q	bS��}S�ހ�8����~5��fY�� Z��kM-��҉LC�Bb���l�� @Q��@��ܛh�M��i�&bΤ�ǷƧǝ��]׬�GE�ԕ��}K���k�BЏ�T]�sXlb ]�j�д?N��������]�8�6A�+������yp>
;�IC��F��m�g	\���D��g��Y;\����� ��s�*��Oa4K)F���K����=i�B�����m������F,Bu��oIR�X�LfCp���tje˛Hep�B�,�O%�7y3��_2��8�����H��6��L�( �2%�
���f�O[����U���y�)��23�� ���h�;b ��7��ǻ�!��'arL��V�W�\�zoP�5ڦ�G3�+!�z76�:��gMD���	�`:zJ~t��/"��Hj���>�7������j5��y�����+���B�_�J$��F�`w�*��&���,��؋��#�x|��u�?[H��fCD���������5N��ڊS���!?-<�B��GvE�`�|��[��)�6Xc܁�$�UV�08WCj|�-e�g��k����O6Θ�R���v��ˋ�k/����"r,�='Af�ü��%Rx�=	Щ��X�̗tT�X��p��xu褋?�r�O���$�~��J]�W�_w��Iȴ�����v�0��H9`�߾uB��%~�BO>�ÃQf�0�A�;:��6h$ò?�S���0G��DJ�w���Z�$T�7bI�76���v�
kT~e��Njv�N���
�<Xz�Hq������gq@����6�V������p�����]���;� ��w��}�le,ϳ��2A_��*@>A祣���Y7��u~�OѦ�����U$��M� n��r�U�1z2A���If�׫�/���#�Q-����JZZˤ��8�}�F�2��T'&(��T�n��4���/�a��1��Ȋ�I��e���巫�10
�ЋO `=M�5�ۣ[n�	Ԡp��0⁤�Z=�J/�H�1M���tc+�)���UbW{�Ix�%�����N$�Qr��X���0X;Щ��&d�q勇���*�F�Yາ���5��=
*�3���'َ�q⢀�t�t��ӂ���B�����K�t�h@n�n���?O!%����Л�#��o#B�&�/��QN��F�U�m�ſ%I*I���s� "z�AX�>Pm���)�jc_�ɢ�V+���܊��:_�Fc��+r��]0��L�n��S0�R��RW[3� �	�'A��bֈ��{aX�N�\�V���Atg�G�R��qV;ꭚ�z+,A�Vb��{��UP���TK��ZU[�2�
p�v�B��G`t�4X��F����i��Ĳ%��/���v�-�m?� 5��o&�(�	�!��C'����Dg!-��I��HJ��O��*��k��-�#�n���o��}��O������e~:|�)��:I@7+*����z����Y�q�3��.k�p�b����H8�P�i��� +t�J�O���L�@ﺸ_�!]P��z��Z�$vV�����ī-����Bp�"��]M���ӻS�zi�y>+;��CCOp���W�c<o(�D�f~�o��f�;.U��{}���H��[V)��U��$c�6�{�&��9��2t�<�N6�_��5o�w�3c�Z��#I����͠��,T��~��Z��n��8�s���[�B,�'�5�6eҲ���C��kj]���+fǏ�>AA�>�Z[�G���|
��C�������I�GZ��:Z]lup���Pz�쉡�F���#La��(T����E��E��U<��� �sكw'�ɡ�P��P�v����I󮔴l"hU�����z?���X�O$E�=I��
l�Η���m��ȏLW�tPCu��
�Ks����	������:��3���;ff8��:�t�kg�\�APK��	 >�J���#D�'���kfE��xu5#���?L�������|�4�B�V�ƈfA�ŁҘI˳�+�1e�o�%���)+�7/��Uv����"�I�6����p�'G���&{.r���~B�|4����Et4Jzn���_җݩ�2�^E(ߙV^*M�d�����^S}i AA;�z�! ��{#,}��=]�/�?�F�;Ͷ�z���:a��m��t���+����O]�q�}Z_�	��A��`b��V�c��E���{��Kjk/џ����DjZ�%
����e���ٖ�qH�3��
pvX�K�tk谞���&�D����q��sf8:_]$�3�� n+���K6ڛ;	ƝAW;�֍��нr����'���9���B��U��O�U�E*���Uq�j�����wu��� Y�����V�$G=�PRa*�;�o��{�A/��k���R:���L`�n�Y	��j��ծ�V�N�/v�a��S�S(��3�	���'��QG|?��*��cD��2�م�� VP5�� �k�Dc�Q�qbq>�H⣵�_/�������v޹��ƾ�:���6���� {�φii������, ^&��'�?�|4��S�&هS �}�f҈n��E�~���ew��ݵ�`	���}"e���<,+Pi1�,���pݜ�����(8��6/�(<ZÿkhM�-��_�����ʟ�}�ֶm�8E ?1�1_̛~R�C�����9fʖ֥ꤌ���4Z�(����!N�H��7w7c29;.�vC[��p#s��FY�^^8A�+���156��bc���ٵ�U�.?J�}K��'_	$��̙�B�����P�~.��o��ҵ������Ѣ^Z�ضYg�)+8�T��|��?G�߾J��3a�Pm}ưV�S�:�a��'�JHi�m,�}�����L��$����Ǫ�-8���7��A�e��R@�h�SA1�
;���S���oWNX+;���4�"��P9�X�N2��������p����
��|�O�����%�=�ٌ� Ud�aI3��,��\��2x��H�p}	�����xʬPcw}�]E�G���Y�\���66;��� %��B���r �l�[@7q3D8�SSCmz8����W������;�E-k�!��m���~���g���];?r��[�P���vD�a^,		�	�xO =��Ԇ\rM��'u�Į�jm�ZJ�N���t�R|���Q��#�g=3��� �w�..�~`��Fy��c��C~b���*��)�ߓi�b���mZ�>y�1?$\�2�z��tȳ�0���������
֋��P�K5>̆d΂Sw['c�K�x�V:����;�un�4��P��q�J�E�O���t�5Ȑ�k�,��� ��M���o��_�'��q�eHT|��RZ��:��e�)��Q�gw��6����I�N�Pm"k�����Pr����J�.�=Q�[�R����,�h��%��� �`~ti�Q�,����f��� S?�"T"�	�q����԰����Q{9�G�C3�?r3^�Y��m6�����u�@v��X6��an>S�x���&��~�[�X�9�a"[��,J3A��"��D8�Z.�;sm�X�ޯn�����!7߅��q���&��U���1����iݯ����GU��>n�iDP��D�JyiO���Ҍ�b8�qg*b�j�#���D�뵁eO��u鋂bN�G�(�ȍ�����Y8�����	�<�A�7\�/$��Z)f�N;��?g�Ƭ������� ��~�R�Jמ��C5m�����|��%#���(@\�x�7c%s��4�;���#��^D4Ws���dT��/b�I�"��>*o_8�D厚tٍ�å�s�N�^'ydZ��~�m��k��_�]��9�&4R���r�;aǽ��J��*Pi�� n؅��س���q�k���Z��t~f�8���+��#����x84�L�� �X����7�3�mxt�zL�sH�;�/���Ӂ�.%L�D��ؚ���]%�g,7#	�n����~뚽��1�lA����G8�h4b���#���Y�"�|�O�䑠��������[���s�����zB������{�=��<�e����O ���0ܾ���
�h��(R.x�E�d祩�k��@��JT����ϴhNX�(ǀP�^��i�a���Q�C��?�a�jX�H�Z���&S����P�5@X�0vt���cj\�uO2��y| sP�D�E��XU_��8� }tp޽��EE��#��r&+K>� �'��"ĥ�3]��x�{m*�����g�I%1�Vsoݴ�)%��1-dI�Ȃ, Z���$خΨ�ȍ��2<���3Oڐ��e-���nd�5�N�42��t�I�����|�&��0�����΍[�eʫ����9x:Tv&���~����:y<�/�_K�S�������z��u�g����0��;ڞ��1"W�k:�z��w&YO�������=}��CN�뉦�:G^N+˿-@��v����|�
�A�`��6�J��$݌(R��}��=wl�!��}�A\`>V�%�Y�M�~E��RPҶ�h9�q��'�_m��Z�n�\����)��;�����'�Q� ����2�.��FɅ��b���������c���9
/�oJ�ߟ*�#>pԤ�:S� ��ҡ���?ެp�?�Ԏ�s��j����r�2��(�%��Ǡ`}8��\�>�}!�kC�lYsxv"s�I�3i�غ���u!mr�VC���3D3%�L��t��M�D܎t��������W�"0HP&��q��W�6���Z���;z�����R�@xBӝ�nt�أ�棑�i~%	��Rޅ/���^��h��SI�'��ET���w�Zo�P)(�|	���J�{`�)'�i��b[�d&:=���I�q�0N�qB8:Ny@�`�bZMy���W�K��;e�ė!�b6˲��vq�n�{��Z��Ɛ�AR6�����b�ꦭj����MT�oQ�g�IaI?�z��+�K���,G�?�$�Uc��f�VX����� �@��<�KR��Gq8��~�P�'C���H�B�g���QU�!u\�g�Y�M$B+�V�����][Z��������+=��k��|_��j��*����{�Gn��*���A
��n��HG����+�Sp#C��k@Jձ��Q��:��:��O��4���TJ�wE��7�5FH�<�����:�L�a��j��YL��]�M"�����ܢ��)�N��v<�5Q����4� 4o��U O�wJۋv�#'�`g��v� !ĸ
��g���uF�����P��C�(�̎�)��^���x:�а ��Aq6��f�(!ǀJr����,
��xSV��t��ôjϋr�ĉ=�_�=�[�#�"D�ZR���s���+��w5@��sʀOL�vń������f�*�q�D|J�I�s�v��\攎��&t�<�cN�N�,R��TR�H�܉��[����K�\;Ҁ�_*��{U9����a� x��sc�ٲ���F����,o��i�O�N���c֚��N���a���ޭ��x1��̆�-�/��?v��N-��A��n!��]���ۆm��'h �D�_��8`�l=���ؓǋ+:�Ya�EXڅ�
�?p�ӷP�#���)��'ՙ3��+���������9Q& �:�A�LS�ٔ  lu��1F?�ߎ�W�qe�｝Gt��0=EE�3�����K��z�Q��������lG�F�jS\��S�̽d��g�NqD'��1����-\�tj!A�C��;D�X1�&���5hZ��]ꦴ�
�i�g` 4�$l�=k�e!wbkf~R�zA��X�w}mC�'�~V��O��K	��������W�T�t(�Z��L�]:Z��>�_c��ќe��+�.\� ��b��^�E�iK�P̨��рUˢz,2��<O��P#��I�Ҹ-cqU�	h0�7Q����/�y�]�N ��-�a�߬D� ����M�2�*Y�zg���K�
At"ƺ>�DǺ%#W�;D� 2Z�!<;x��A$$#ɕ8#�Үk�\�e������f���}o�Zc�����y�9.�Ҵ��\O�QE��3ɧ�� �k�众 �yh#	�=_CL���=��wf
�K��3�R�`��H��EW~���ҿaQP�z$�N1M�]���3��z�����(? �:�`ۮ���:��$�Ix8�<7�;���.<C�ڃ�I�^���{k�E>+���f �邲OgKh��WH%�� �w��"��9�ϲ��ɔL��s`&Cc�(w<����	u���ο�y�Lz0�l^Fש�95�7�_"�����ǀ-�+p�y�*J���"���#���pnL
�&��V)M���R�Y)������#mU=��c.�jg�_}�HuuE�k���P���t���R�`n��8�YQ�x���/[N��C^ril�^�F����rt(\�*خf@P]L�(�=�)��D��u��m�
Q���s����=d��.��r1<F	9K���C�����mA�\'�K�Ϊ�јs-������2�YB��J�H�\��@t�6��O���4����v�l��An����j��ءz�� �B�t^@ ^w��$U-��0B�H���wՇ[fl�ޤ�в��-�'CAo]+TJ	�T�p�o>�5�tX��Tj[f�M�^0u�9� ,��b�$:UN�J��p�OI��U���"�����"M\}��ѓ(yGw�x��i8i��rَ���rI=��������[����="'�H��J� �i� ���Xf�����P�\M}?�,�Pu;���q���F�o����ݡ�r�̋!�������KZ�%�.FQ���R#�[ ��@����!wQu���
 á��jG��+����WF�Y�}hH��{WI�;T㇁qFD����CFT��/�}:�����&�������0#??D `��;��?����8�4�w�Z:O��٧�E��aJ��f2�x�eR�r]��k��;=ѹX�f���L�;bF<�l�.o���w�ٜ���996����2��4�n�F�
�u�#�;��X/bB���q��]�-�!f	W�zd$��!�L��' ����F��P��&}��Oً�6D� �͠�)6 L
pF\��G�בn���(bS�1������la�+?^몲sՄ��Q y�Uٳ��&�V3������n%���2�����)D�5�Jz�x2� �}$�ǻ�A�s`�Z֦Bo�B� ��`�� �Q����~-�iL{t&��:deW}J�@����'_G_t���F�9ޚ�*%��]�[+���ߑ��`Ư���u:lu
���'&4�����1�P����9�L��4��a5��0g�����Z(��ﻶmQ��)����o�
���� ��p�̑�N�������lc�4a*
{�RT돐���)�6$t6�s��d��s� ����&6h�"��ǎ&XtO���/ʕ�����7l/�q�4
�5�	C^����ݩ�W/�?�߯X���X���)��X[��.C�]&�B�b���)ֲ�>��k��fmg+�5	�' 4~�(Չ�ۊtߒ��n�R���A(z8���r�G�����B�6^�:DďRS)OHs��2�%	�����f�����`Q�2��$8��E�+����y�~e�
Z��M&i@�j89���Q�#�������[���aqƘ޽v��M�sH����V�>�j��B0�ǔENU��me��T�P�����T�!�,H1�����T;�y4|<4�»�hY�ci���,�@3�Q�;��8&�׵�Iö(^��b�ٳ����:�g�y��0��_4-N,ك�t���|����mY]�
�Z��2x>3Xa�W^����/��ɹ긽{ox�*�p>�T�M����R5�)����_��>�ag�3�y��@y�+#�F���IRf��_g(���0�i��F��{����ʬ��!��|��K���m��"�: 7�����X�<�riM�$�cdz��p��y��? ���-Lv`�ޣ@LEYJ��W$N��y�$�5�P6������+�b���W!�����[ry� �z��*��7@���C+��
����ʸ;�q4���)1�b��}�n�7�ڲ�� ,3�ݤ�M��������jp�5|��T3q��:�׸k��L�4!�U �~��p���5v�H�+%�aQ�[J�{5��Jh3��w;|v�1�E��/��K������C�l�%+iq��U�	�Cac�i�0���A�E"Z�z���3W�V�ț�-��Z@M����P��7O�r��J�g��e���)�'3O2T6{zB�"�-�u�Ǆ��	q��_3
`�Wㄧn�$MN���j?z��{��@lل�ry#	\�D��j�D�wQ?�0TK��+8�{^q�ȍ��1�e�����9;&�e��o�����ӫt=<s��0e䃚�|��7�����uF�kvc3�y���G��Q�fR�ZF	v����o?i�D$�E�Ų�����T��?z`�3���@��s����v,O(?vݻ�l����e�Ƞ��H�
0LuG�~�S�nd � �>&5�Z�`��t�c򓣃8o��{�)P�V[c1���|%��p�&���mQ�[�F|5�\�|e�NTX#�Cxg�7cŚ���]CՀ�O4O����W�X́�_��A�Fz�S��a q���V�o��`r�xO1|ݑ 47Z,��lrbbq��p:�2���Ľ\ L-hUJ��S1#�d0���P��Zt2�qٷ��V#c�uN��UJ�h��bc0�|��ii��M���os��Q9���C
�	���̴~�;sЮd�1C�>]��¥*�E��G���ɐV�m��W@1�&�
?��ٳ�D�v�M��a������8��tn��Xx>���+�蛤s#$��$+l	\���M=t"���%/&%��������%bH�zt���T�C�TgM�7��D����+'�/��)=븟69Fm��F�V���f�\��t�Ս�����a?}��f����x!���R��P��d{@�H[�t������Ҟs7،.F�eGH��,���#��R�谑%�.:?k���?��&n�(Q�֚�W�0b�Bl#;�T��^�?Pߍm9�^��nC�!X��wd�����.�Yr��z���5�C�g���
U�c�`�h�A�ư��H��EoB'�#(�(H~��(����E�?���R�b㮓���:$
���̢���O������_��d��m�y1��1��!?�Y��C
C7���������&�6��=����;��dyep�#rch7jL#k��������S�T�s�}`��T�]�{�DC<�&��.�j:Z�,~>��Z!�w~�� T�����}I�F��{Xc��6'��.KS�r@��9� �@�� �Et}��

���blW����85�'�}��r#=�[[�vb��xk#4��3�� ���P��9���� .b���t7i]��ub�B��]�F��[iPIQrV���@&C�p���TL���@�����%>��th����p�P)�}����,�>��v�CX(u������,,ύ�V�Kh49sT����̝ĩmH����61�St��%�b�<X���
��8�K���z�����]I��a��3���v������p}��p$���������i�e`0g/j�[�Ψ���kh�P
R���"BL�����۴��(��0kh��"��~�d��ꅢ+(�;<M�Xh�/c�ȃ5�̇��B]�h�qT�K@5�u�_�g�}�8���w�z�i%^= �V�fp7[s�ڱC��7{\��U< 돌N�B��Ww&)�v�,�J�X�c]7�k���A���w�����"�AQ��ZSr�$J�J�)��+���"?�.\t��"Rٟ��o2q=z���7����΃���+��Q�n������}gWq�l��}��V�Y�y��ø��	��Y82�Q�l��p{��\�ꐭ)8�i���S��1�������1=���=��{?c+O ���LҀ��Y����} 6���;UAx8�q�j�^�<u��e�6iΒN�Ɯ~)�-`��D����d:m�*lB�^#^p2��F��H����TE=���j��׻�"4S��jR�K�F�8"Ujؙ艼���b�X%���,�=����R0q�BP�Jq�G�9j��:T)����9>UU��xȶgZ��vQZ��rT* >ր< ~r;��.���T��h⏖w�ȳ<���ĳE�\ �]l&�<Y'����,�"�����A���Ak��1��ږo�l�"  [����1r��K0Mgmא��t
F9,YN(>	�nJE�j�c�y�<�l�Ty*��B*�5'!��/23���)�t�D/ �	�?��Ȅ� �.�����u�[��r�i�?F(@'�}�� X��h�������\���k�ÎJإOߴ�������sT�`��ʷ���ET������r�<J1�ū,�����T�խ-���K����T2���5GXN�ljⲫ𕫰i2��uH3���
�|��~9#R-�^J@�Z�CՈ;ɍF+a���(%Yͪ�o(GG�����]���زҢ�ǡ��� ��*����ȡƽra�0�a������B3�4�.G��e�&�)�`���4BI�Na�Ėc�^�'�+]�1����*H�fMc�H��C��I��J��d��&bjCbƐݣyX��AW�J&�Z^�@��HM�O�(�h�%̧P
SMӐ$Rw��|X��H(�
g0e�Sf��I�R1�5�m��~N �c��G�m֜%�S#����[�|�KpznWH���g��A?J�2F�>�]���3�E1�o��ܑ}J�{L`+���)v7}�k6�w|�g�/���j:�|�=k{�w4�՟�Q8�EW�+���O���.<�+B���wgD��+2��҇�)��?^b}n�W�C��c
$�>�o��1%�֦�X�����D��wK@	(k]�"��������
G�5+��CF~A����
������4
��u�tƝ8}���Æڠ��+L�(<arX.�%̔��7���Ù�Iބ*w��2�#��0ʱ�g��js�W�AK'�Q1����)�cj���-��Rx�6�
��l;��U��MYI0Je2||PT���w
O�S�ےv��5*��*�
N�i���]ֻ�J�8',�ҧ}m�'�wհw6��BO�����?���&���q������{���קa�9਋Q�t���ź\��O_0�Dk��,Fg���P�����R���Ou�L�'T�� ˕x&?˴��\h��Ti^Z��#91��\���4��� ��sQZ{�!��m$�G-�Hʙ���,����9��9N�c��{l�iq\�����Q�b(5k��z�N&T�����|�(�����I>	�������*r�ǝ�u�oFV�ju���K�1�&��v��u�)�r���I��g6,���M�/Hfb�/H3,Ó��Vʌ3yp7BO��b�s���-n�2<����K\a��`s4��bb'�C�L[���B�
��=��,������nxm:g�n_ <9PW�^�/��.�B1Lc��4�G{�3�j�аS��dR�^=e���'v���v�vR+���sv�_'�����G�3��_���.w��&�S;��	���OXZL�'�ڗj?�LIG/4��x����D��fdE3�c��ۈ�5���!H�d�~�Ze��R�(�W�	?~��IPo|	�g)@q�k+�3L����SP![{m��������#"�忥�Ƹ�ܕ�`d��m���v滌8ܳQ��� ����s�,8�>�-t8�i+������l>�����ӽ��'O8�VF'�����t�����Dm��n�a7ڲΥ4Q�j��!hL�8���q�R�K�pӶ*_�24d�$n���p3]���Z�Po^�?5N�����?�}B1�s�����>�#z~xM?7@�c�ɧ���k�)&����N��MC�L�X2x�h��!ԛ�b=�q��>G,�P͛��f���CSq����ċ�@f&l�ֱA�����.������҄�V�ֹ�~H�w�7�Gg=/���d�����Ν�����?�%^��m�<�m��E�J��c.r.�	���}|�����l��!�#Vy��~ >���/��~`%�:%@�]��8ưΞO��sT+�2ICf,K�TT��_%Y����� ��E�����_�9���:L���Q��!������قzl+
�����ZZ��y�`�7��V-��T,�ԉ9}��ܽ?��$ڱ!|��#Q�u�s��N�Fb�~9�S2P�E�⼔2���#�a5���	 �H3��c�y9�!Wd�7+cl���
,JfE�8��	�l�u���1&iÙ�aj�cH��>�L�t���W���I�+g�\�Lݯ��X��q��c���vr��3��^<�����p��'��gr|�*P�L8P�ϰ�y5�~�icѴ�ؘ�%���h��:<���O�.E�����e�1�!�u��އ�[��^@�Rs����V��C����t�2	f=� ��a�)�M��P�v��R����gj���������m�|����t�ʆ�G�yY����{npX����KX�5����p���3'ݜ	b���(�|��j��=;����y�l:eL�pٛ�;6�ǖX#��G���8\����aC�*9>L	�T_�h�` �����K.v+�ֶiڮ�=YL���љ��!�%h昈NǣN���B��{�T��c�ƣ���1.�*3���!����%=�c-E<u��*b���iЌ�f���y;����SE8� �1$����C�:V��P�����a�y>��c�	�ѧ���qU��GS6�J��lr�|v�����ӭ���_6>��#���X�0q�$��K9=P,�������;u�Q��"o#U>�mB���.vV(m>����aC�1�B5ګ�Wހߨ���)uF��Y�� ��=�=��4� ����洪�Z�Β�x3_[��{�1���TJ��a3DlT�������f���ހ5����g��[JO��>[ݍ-%����O_T�R�c- G��'? ��zZ�ȔrN����ڊ�$��z�Y�2\R�5�|N�Y��l�t��l�/��W]u���۫��{-����7N��OB��5K����a8b�3?����%z ��y��?�\a�]��E�a�Qq��$��&i�8W-n*� x���l��b�G�ꀰi��$��ྙl�u�4;[/���ʈ�%���(~f"����C�Rc��Q�=#���]�]!��W�!����h[��ܭ�������s ,B���}$�š׃ʺ�q|n��w~�*5<��G�8D����ע�8T�j�Um���2 Q��M�A��� .�{ӧS��_�(��2�'���7fI���h��Y��+�m�S
��s�9�Y1I^X���V�ݾx
�)y���c���MD���Rq�@/q`)*�I�ˎS.o�T� �f��R4��R�n�GF	q���U_j���q:S>N�����J7=������-��K3��7�S���D�L�;�}bP� ���UE�*��)����,F��F��^tHc�1�����ּ,5�b(�
?P�k�%Y�KHY�Rcp]��5�q�n�R�x��<�����(�_����M�@te�sx���#㿁A[j�v���*���u�e��%��q��ty�X!�����h��1��8��Pہd´�:`�ؑ�l �.���V~ǒ0C��T'X�TVWw�I�F����Z��U8��֏V���hQ�S��� 7}��+�
��������WC1����MN黗s��=᧥��yDb���[
��m�{�w��&���H���0=e�vA#s���L ��>���,\���*�;�f�K�K�xV_��`���[B�J�����z�G�C4á���F����]���r���RG�V��v��_���qp���)�H�U���(���e�ǧ{�.0
Gx4(���1&�������z���3�Y;͠�VATr-�\�b�>tm��:�+������4gj�2��\��!�u=D�@�G��w���F�`���7ֽ"�d=�O�-!����$���u�s>��x�G�}��V��Th ���m�!Ј�5����׏��
��ړ{�� ����,�ȽϥiV��t؀�g��E�)�m�~}l\5��c[YC��G�����j�NFnv�.{Ag�2d����pT�3)�{9�Z���!��i�1;~���+��|ƶn"�*P38sw�L"v �A����|ml;������k����-^�����)���Gg�+�n��jG|%>#�c�2�o޳�ϯ�s���i���V)�iܹ��݂
*h0g���RZ�oϒ��;\��z#-�~���؇J��O�R�N�4u�rs�b'��k���[_�xu�ұ �-]k}�]�TW�@Y�UE���Za�9�]Ga^�4�\�gԽh�f���T-x��0g��K1������D�ź(�2j=��BU{��*����oX���ʂS"
Y(�vK��M�2V�i`DG�Ű�-28�)����8:�u�3c�=���#[�v�j薩���AZ���{�c,� �ڇ;q'�Z��n#�*}Հ.�g~���	�`p2l������ظ���@�<xZ=(e�2��*{���%�����W͉�����?�B
���.O�5�++T��Ji���t)�4�V~�0K�Y�n�Z�y.
�aIy��^��a0�ً���e�TD��һ]���Jƀ�X e:��K�?!q?نt��Oy��{e�X��_�k���X��5ޥ!�Ba���L�:#��i��)���<����LqRŎ�5�Ѽ��$��R�ߏOK�3)C�T�Y?üu�#�����V�
��e���s��?��Z@���MF�����
'��O��q�`�K�!��[��T$爵j�x`Ir����������=�3��'���3�g���=����~k}Cܳv�_��kG�V{+v�񎉃�F	�$B�f���5�^_POAÎI����.�H��xָ�k@߳���^�{[^�㘏�����I�f7�sx�(��a.�L���`����A��c�������?GO��������Kc R� �֣O4����2L�h���:A72�UZ�P��+M���7�AEz�:;:~{��{�e�W�''f@�����ޖ�lWp��u����}�o�#�ņ���vw1�W���4���w8LJ:��j]T�a�6;�~��7�����t��"�D�Rx�Ii�Ak\g�O�TtJ$b��x��c�.�}�Mc�6M'���<X�@��TR����S�rSDBGQ�V��,ź�4L6g�xT�v��ϯq*�tnR)t<6<N�����;H�W��ϥ�r?L�6�m��G��a??��S���R��[�QD�l��Ht�Y`Hl���xZP���?^=��)� ɠ�_��!�y���L�q�1�VQu6�\&�_��|�dy�Qy���K m��C�5��˸t2�B�̍WlIP�ٗ�y3A���quUҺ��/!��Q���3q�Bm"E��U.7��@�C��E9��!y���&�;�����F�$�Q1�*G��
B�uj2~����8ڧz�!Su�$L례ێS�ot����;n'��@���}o�;*H����R/A2����P�C�f��hf���2�ʒ8��ÕɁ�*4E����HI��+ܚt��1%|�3|�g:u�����3U�%�앚Z�߿ڕ���@�a�(��?u�b\Lh���ɵ0(c_fA�ᙊ"&�w�ehΞ� 	�?3X(	�_�L�����?�#(e��5��N��?r���#:igE���nwq��`ΆN���� C��$��-�ˆE���d��<�L�����]��j�d���$�� ~�� 	Z�H������(6�J�9S�ncW_���6L�7L�6��%s��V�@vv�͝E 3�C���9�������縆��#S"���4����:��t�Wm�
�s"k9���4��%ՀXq��C�=x-�C�%�O��.�\�:�^�O�LD�2Α���w���rݝ����ß�;R���d����?��L���ԇ��u���A=��y�T��`p�ƱW�E'.���}�ÁB��w�P�h{��e3x⣮8�w����&�eDw�h�e��En㯞��������0��o�y�)&��`.�]픲{�}k׵m�Zou��e8����]WK
9q��k�tE�[;��l���y��AI��=��.�"F?�F��lj�Bs�w��[A#��g�U�0p�Zv�@Ң@譕��/Jb��,_���In�V.4��$c�,��/H�c'򬅽U&o~�3���;d�*iMlu�^���;�gޜ3��l}�&	��Bv��4��Ӯ�&WɁ1#4�u����Cl�ҝ�s��n�Ek��M#˫��� Z, |�i�tgRg&���� ��旛k�i�4/C���w�i,����,�+5�% k��9�!�7��Ca�R������c�*܎�RC*�]K:�[�� �YTu��¢��~D�,�u�6>^�f�W�C�u���GV�I����@��5�q������v�N��^|;���S�1.��dO�p�J�gR�ܷr�M�g�)2��ोi �j}P9�
���|U&+�~ۅý�W���^��7C�/uHJ͐��"!��$���%����kv����R97)#���T�=4���9�og:��3�kj���B�x3${�P�z0�>q��RʪBuJ�
M&�i�1�-U>=��3�mZ� �.�	��V�i��R�zd4)���#2�-�����i��5��Ǐ��|^�~p*�3M�R���/�K=��R��Ъ&^��&�:TDNw2������� (��ԋ"D*3�sf��[�ǳ����tpC�|:�w�d{����<Y�ͮu�\{!X����jb~���e�ҽ�>�1WV~��7��8`��6]l6;��b�8+�*���VG������ᢎsN�j�K|Wo�7I��cY������1<.�X��g\�-}@6���LJ�#6<�x6(-P��M�@/���V>�\
��_sE���Ӏ
4`�V~�iρȶ�t�� �c�ì�AG֙������E�|qO�X~�+��:�1=N �A!~��Okx՚�����'{���g�K-0��;k��eN~�w��R��{��B�<;>ea�s��U4dy�_�r�'VVh��?���Ah]�<5�4>�y���t4ϼ���u޿zPdDU�����n���Z�[�$����2Ȏf����|����~3�j�og�NG�W0�(�{"&P~�Ne��g�����D�U��e}q�))�
�Z�y�>PХ�d@�ݕ�{q7q�/_>��zͨ<�o�U:���$�cĆ��t�ys����+��z���F����'���7��E��*��@\�����B���6�6��(o�f"�H%��u�p�i7�k�{�����I�ěb��JU���/9�۵�帤:߿D�Bx�=|{&j�e�{؁�#*������逭`\;���
"3�^�Ki�8�%�B'S6�U:�l��� O�1!+c���� ����f
ݶ$K��:��*��KGOS��>�����6�o�/�]�� ��FŁ���C��n -C��|��h��a��=0�b��$L����v0÷�5�()a9y{��ۓ���w+�D�s���-��#(R����=�
�.Kd��ߏN|�~��CA���u��/�g��O��V�+(�����$"悬�4� <^L�#��V��Ba���-�M��:vX'6#���[�x�]N�pl�#�7{q�o���k���
X�]7"�}u}���p��N�x�#��	Ґ@�G��( ��{����UWVe6���#��2�P0*G:ю��k���gn���k(���is�Eހ T#��K�@������+���X <%�j�=��	�^����m��@Rթ%������)Lo'�\�^k{Lh���ͦ_ST��X�Ѵ�`��d���#B�L����G������`ml��2�*�
�c��P�i�b��e�h�Կ��+|<�Xh5�|V�D/��䘗,��3�+�@{��-��+hxz�$�����`�X!<�#�Q�svj"��euČ`�K~��p6b�ť����O���kg/v�\Dh��I����!H<6���U5���<Ŝ=��p�Bf��G�B�� ��&N�dę�䗠�L�G�,���t"=W�J&���m6bu|��پ�*���g��G#����֯E�à�b����?�<��NL�ֽ�[\\�xQ-�82��]a��0"4� �8>��(g��2w.�nV�5����� �3�*#�6�&T�O+��G��O�!��#c!(�3��ON�i�u�t�,]J\l�>x���8�����
�z�k����O�'�U͎u�|X�}���K���h�mO������'^�D�Z�3ת��O�(��9�[߅��~�;�&*�ZC��@;�l�;Y�t�r�?X~�%�z(:����kx�`_	-l��ƿ��yNyC���Qa^�g��hH�?XL�Q}�q0{��pQR���D��Čq�5{2���k�Zr�����՘�o�K�+�g�A�1=�b*�SԎ3�X|nR%���QQ�y���|Y�a
�J�� k��"Q��al���X��	 ��5��-�����=K "%�����lN�s ő7���v�����Te7�6��;g�e�S܇�c��u��ҡ��1E��� ��+<���խ&�6@�V&	/�t�As`�a%/���٬Մ�G�2�2��.��?�����w�KRF�TU����'��2����v��Fս��= 9�hz��G�-��h�;&�1�1MM�ݔR�{����Ǳ�ΏN�Z��m9��F/����.P���pM F]��������H|��ok?�+���2�_/I�<��p_T5P<nmpƀ�[rN|����B��)Z��T��|�G��k7s��u�ifnV/6�kY�G]�ZDL�R9H��������-$��e��~9���a/�r>;oq���W� �-�r�P��P�/R�ȭ�;p#O��X��h�rq[� �?��^Pϒ|��~���P�;��a�`8C�dh��򲭙�m�e׊�"�3���y�� w �}��D�$Y�w8L3���»�'d�%�&/�?��w�Ө�)�X����f��dl���.@G�!��TVk��Gu�a������%��َ��z��
ł?�1֋R��G�R�:�?�X��}^�gn�S�b�(|��eǽ�Po���{û]I�|j���)J9\ ��UL�.�{���9
�+�~�%HپƸyi8���9��ϱ�����bu�?���v@6nu�X�z�?`�ʲ����Z���?����NH(EH:ᱞ��D�����s�ݱ�����˨O���c�����E�e���.� ���C�C:�So��Q��[�j�sg�\Q��Ø+8��NܨJ�G�5�-G�uy���L��ʝ� P'�"�f�Ͻ�p=���t��M�^�]�Q�Dt?�M������8�L��U��x�m��]����A�[���(�lQ��?�h�UMiF:޿N��:�ِ��
��;�u�8gG���6j�>����w�#�c�pe������GC���y��W kW�-�ux��ˇp�-h�EU H{8`(7��f�{��3�ݯ4]��A��O#(�j�R5�d�6ʙ����(��T���������T�L��/8�V����ρ����M�3��}`�[d��s��-¦�?r&숺Q�W��wW�k�¯�Ò�k]��\�����#����]��E�ȸ�*�/�ٸ4s��I9o셽ifB����	5\{�)����x�R	�b�}-�Y���`��U%w�R�o���oW�)2/wf��G��K�TOP*� �!�f���L���/LʍԬ�B�9</[)��&���Ė��ηüw�_���F�X`�O��}�t�~��������~s��n��m:��<0�ٚL�,�����֓�T��>{;�b��D,R\n�#��Aor�^�0$/�` ���h�)�1�n�RG�6�J�z��c���D�(�a��74���jƘ
۷�/D>5-����ʿ�jx�_�jd�t��wvp����s?o$�Q��Z�Q�c�%^<�=K � �˜���e�d|@�<{����9�ê3ݿ���]��NL��'&l'�/@��e<q�e�ũf*7#7�Q��=�
�<�u�hN{~����ᑨ��f`�Iy��z����u5\6�� �Pa�;��2�m/����,��迚����h��Υ���V��������v�dK��&���3�-򇏟�����ZQ�gZ�R-��U׊�S<蚱��ȫ�(�I��/���gT��PV�2ҡ��f����p�]�n'@]�T�8b�?�����m��UTm�����4a�M�<qf {8jO�,ޢ�6~b>���h���^�|u��~�m�z�d��{4�x��+hQ��\�/s�s@���Q� �ż6-g ��͞xw(ߺ�[#�������<2�����d�*�FU��p�{ �qjG�#�y�T�ˁ����F�H$:������⹉v#ۖ!��-f�M&KB kqUq�		�&�ޡ����xŁ�{�0�J�h�����b	�W������҇��>|d�J}k��I��|�|ޕI"[D�q�i�sܗ G=*~d�MAn�L���T������+�=�'Y���4��g2���3_^�d���3��kF��r������{	'�ti�py�ٳ����8��>���}��˝�N^�8[C�Ƃ�8�嘃�8B��ȟ���E�^�����Zj�zA��ģ�¶G�k^����*�Zx�8!�_�}�%-���(�M;� �� �(�� x��I��c��ICl�X�A ���j�k��O�&N{�G©�n^�勺�m�(�g�ー)���4����j�t��c�X<���d�y灇|��: [6�Ei$��O_����>�bց�Z3-�1�-m��,N��u��w�6�8�f��u�����xIavUYۡ]��LC��w�������)W�|�����C��>!��a�ou,r;Z��B�mR4Q]1bdJB��/]8o.�jQ+�v:X��A�����3��bf0~TG�����§��L�Q=����`�.��F�;���@{��T����5�ʱ,�|e��Q��R�lȼ������{s?88~
 �Jy�E��ོ��u�@|��"�>Ohk6���Y�dz�D���~k�E���>?�H�:*JV@��@|p����OVQx(5X�2K>��ʴ=���~\*YQ�� �1������XF��������`����`�
ר���
H�(B���>�Sz
��HZ�#x+tl����@�\m<홳��s��p��m����.�& TB:}��������W�D��p��.�z���i�pIiIZ�~�  	����v������'O� �f��8�$gy��"�t�D��	S���!��,�F����^x�1j0�����|3/S܃Wy+V�p�����*�r�T0���dKH�����3;����,"�4�֝l	I]���?���>F?T�=�-y@����Qn�FH+[s]��!xR�h�/����%�����/�ՓkW�w��q�l9�.t��m�RHMeI�Q�U1.��'_z��/s��k����D�/ɥ���'?��9�)�,A���Q�/����-'	@jP�)��Y�aV��7�C�5G�[��t�����8N]	ݚ��k��VG�o<���KH��B�It>n���^(�XZ�}�'+l�����x.����S�m��:���r�3�l!LG�� ��څ��f\G!T-K��'���^sak�R��?��!{mF���@i��K�X�1V�p�%�ã��y��d[_�V��00\�t��L�2��9y��g'p\kC�΍�a�p�8�����o����	$?�kN^���;� Ԫz�$�����cuu�:���th��9a��#@ï��4�jU0FyC�6�Î;��,�a~�v
���'��麏���T ��%����ȣ:FkeE@��f��8�Ǣ�t/s)&��5?2�7����!� n�F�i1����v9�Ly12&�eDp�Ҡ�R��l�yϦ��d*�zЧ#٫��hX�
\D��pP�M��q���~�un�ߏ{`��d� �C��5Ԫ��N$�n�N�T=���_��<^U���t|U.��!���w�F�f�K���;�M�"��+��V�	���r�=��F<2�+v C/�QT?�&���[�8S�h�����YiЦ,!P�ǎ`�۹�'i{R��,(��,��wY�Bl�e�k�$���_��Li���Ηyj��-�0{/�؊�� %���v5�ZemHh��x:W�wa:V����<|�장�9j��%���S���g��Fn��/k����%Fw��^���ut�ƻʎj���k?l��3$#�^p�� j7jkoPQ��U�w���'أ?B'�S�W�A�m��h�Ar#��`�t��� h���h;c���S���f�"��D� 5 W�{F�-�*�[ݹ�]���_�!��>a�pi�
�b-1�d̸]�䩛|�ҭ⥓�
� %�Mق�7s�r.���j���f	RD�{��%�L���#����xP�@��f!��A��:s].h�/�M%�����UD��p�D��_`�X ��e��4�U`S��b�bS���6n�Q�Sì�j:��i�ǆ��1}:��I�Mܦ~�=�7lݯ�1��0œ@��}��况��� J���>�� $o��S-A��.�e�}[���6��N6_ ��9�#�0�q�:$}v#Q4��$'ϧ���ϱX��D��BuU{>lM\g$�L��T}��eS��:@jeW����4l�
(�q-��{�ڎ{+�d�� �7�)>�,	�F/�͎���ml)9Ͱ�^$m�h�>��߯�/\St��SC��)�����ܯU���n��)���Ig�����C����'�͡zq��O�u'�%,�h���t� �5y������b�`��"ڔ�X�A���Ҧ�o#�<)t��Y ���I�F��T�Q��(�DD����($xF.��Xy��J��k�oY��,����WGdb�
i"��S�q��=�����N>�5<iF������lʝ>�H��Ypp�O�F��:�a��޿���8��;�����ϕ�X����O� ckcM7��ރ�9�j��@�OP7`��kWΞ�C�~�qz���~�J��`H,����__�ɳ\���o�3�)F⨼:|>� ݧ��
Lc5���pNf$�,
���ؙw�I��X������E���Bt���!�;�ˍ�`�|�
�7��`H
��+�����Nca���Q��h
~��I9��%�v�i�m�!���H�#�C��#��scȨ�!��t�ng�DgNCZZ%Uwd�	7w�XW�VKX�o)��8t4��"Bu�(~mm�$��� 9ʨoU��������w��T̡�#��E:*z��~�{)O�I8��!�\�DYʡo9412�YG�Զ�"���������s0�l�����;�*��y��/]dR�N�y@���_�T�����i��Tb�I6����Q5�w�R�I��ī�҅+�g�"P�D呈��n-4툙;�
�����>����JR��W�י�?dO��S*��'e?Ɔ�Nh1�+O�_�j�|�1W�H<Ǯ?�}G-B����UZ����D���g�&��Ϊ���մw�n�6��=�� �fi	��^���54�h�U����rF��Q�skL�)u�5����@X����Ivu�+�v�,_��|)z ̍T�x�G\���-�1,������Y�}8�E�d	���P$;T��R*s������z��ڍ�h�4�~�I4�}���N�f I�!47���X��i_!w:�r*>�v5�]"����tPe{"�)�(���]l~=�@��̏�����ơsŨ�u��N%��XZ�I�h��_Eq�@".%��sY��h\A�[xM=�H�'��]���<�a�V=2���]$y�|=q��֌X�nQk]b�vi�_�V!�-�?B��s�ǒ�L^�at�3ɍ�ѷ��V�%�	a��Y��a@��-�_bS��W���'�X�q�0_��1�l��[� �m}�K�J��A@����QyP���Oي� ���*]���i�po�p�a�nfNھt�U���A+xO9��s�~¾у�v��u�h�ڇî����4�>�bN��GO��BltF��)��$#'��� �� �^�]��g�ų�L�҈gt��r�;����s<���Fj!W�j�EkB	��]^L��$)�B	�"�bs���i�����֋M[����k#B�g��׈��>7D���q��_B*��5w��;
w6&���R$}W��K�o�4�U��`���,���fW&l�Q�t\ ��Sɻf�#�v*��b�AOYj㡻�o�}��uKT��M�ng�@ �4��	��Vf��$yͪ���`�*K�&ǯ64��Y�%��_@vm�Ge3�����������Rr�g�HC����E�������H����	>N�
:j�]�P`�Y��j��K���	F�G��x�̮��))o��wM�����H��:���B�����[�#3��}���d2��{����������%���ڸǤ�!�,�sZA.�"y �dw�$�Z�a�O@3���FMC�7�ϳ��X�I�����L��{/vӱ�<8R�,2�PBlj\	G�șJQ�+��'����@����dg�هX����c�jِ���AtU#�-=�h ���Xޟ���b�{eX�nܦ�7�@�06�����XF҈&?�X)7۽67x�P����ׅ��`��CI������'����s9Ї������9Y"��}���_���N��L9Gh�mIFķ����RO����U,���]C !։u�����a��*q��FY�&�t��=�ˡC{�rm��	/XE�r��DG����>,�ڕ��4��JQ��u��M}��9�:����-��SoJ�P��V�������Ya0k�z���$֙��r\�<'������5��`5C���e4�����I��2�R�Y:=��T��ە��A�J��&Q�]*̵F%Qc4h��Qz}[.dMaΙ�4"~�$H�L��6�{��L�J��8@�$p����� �����6��wMHK)�������z��E/�{TE�����&��ӔQ�~�_JF�-0YO-�$��C/��N��E���t�/��u,�O�O� O#�|m�=�ͱ�����qפa�ȩq�)@2B^ї/x�@���j��_��z�`����E��X�fj�N����h(Gfv� U]6ۂ�\������'�<;=s�@5m�VJ�w7��8�q��A��<Ē�x)��>��`<D�� ���(��i�8���Q���Y5b�!$�UP-Ӻv�)�<4�Ņ�Ӂ��x�%�4q�����X��H!��e�x辡�i	O��F�w�%!���Х���]?�Rg���M��W���si���v�H�p�[�� �E1Ϲ�
q$�c7�%���争�[��U"3�ޕ\����d��Sy��i[������UxD�2�^������o�Y;���R�H��߭�ԶT��y_�iQ	��D&�7�V��#�H[�zT3ٴ���.�e��6N;�r���P*�Z�oj
��Kc7��_M0͞�s�+u���n�C��g���2/hrK�E��>�oh#��Ic�@]\S���"���<�!�H����+���_N�����"C�e�7�v�7˵3J�Te�FV�}=+Qӵ�jp��⪘�� p	A��`E䟜�MJ�$�i��N�v٘�.8O)2YTԕ���z�oP����b����(p�� �ʽ�����,�M�H����N�U�6��(�@�����r�j�>L�+�wr��R.��X(`*����d[�*�^$�yd�'��J9��� �k5s�Z$@��w��P���4)�5}���;"+�-E����**�I��Rmq"��H��僗d㌪�OE߰�#��{h6�Xw;[�j?��]���̛j.J;r�JP��ӞSZ�;�=�cV_��R�Ef=-��;;�}λ,f���c���f1�P�C
�=r(�s-'��^�!�*L�VsrD�9�����	��@���{�9f���f��Z�z�"�!�̄�� ��d�D������J M;��E}w��	�����z3���ح�d�]�9겫�9�snˀ>�q���6�6p�R�jQ�%Lhk�"WH#�Fe���Mė1"����L	O�~df�WYd+���]�]�-Č6!M�힌~�ƣ*���|9hH��||��P��IjX�>���,ņ	*?�q����.��F
�*�&l'�RL����Kg����~n����͈��D�b�+�.�z���ݨ�6DpE��6(�8�c�����Fj̟↎h�U��N��yE�n�$g��Zt>�Lg�����tB���j���s��7̭�?V����	���gw����+di�,��h��q�ڛ�jN�W���.��}�>H#5��e��D�u�Vh�ێٟ������@�ch�0q����>��]�����;d��M�'�u�cE�`��	�^{Փ����x-�����8�Zѡ��-�s�<f�b���a�OsҤ�j���>��{޳,�
{�4���֜ipLNz(c%Z��3��UC_����C|a��.��9)2zGK�����g��!��H���7p~!����{��-�o��n~\<�)+R|ɜ+�3� ���	I�P%��*(������3�`����)��?%��o�1�@
�t&w������ʽ�b�����B$P�X]us^�}�b��6�E┃�~�(n|&���x�I��5;��Lϓ�^��k0�o
�����[�ipw�-`�(�jQ�F��]����I�UN�8T٤��t�I�5��ώ��S�W��RƷ����ѱ�$`A�y��C=A1��c�V�pn�LOv�ʭ�*�w��v���i͖�T�o��L�V��o�'��Y�\L�x�P%{���I�^l!�����f�~�!���.92���>w8GA�]0�}]�����]��h�
���VO���K��f"O��rSUW�x| �Yh��ABFrqe.9�v��,n��=	W���,�H#�*}�4B��?�b���^�	�MQ4G����5�h�TF�t���#C�nR-Q�c6ǖ��2{���fcc���M=>�]�O\خ��o�h�6J������/M)l��_�X�`�����`U��+n�k9����.M���Z-�S.��� �����V��k�t]R�p�0=&=�m������
�P@��zt3jv_-� �����~=&��1�<轨�
5�5�^� �f�Y
bZ"A���A�&�宵��W��C&�J��j,�%V)�����=��ư=��5�2!m!!�9p6�x�!�����}H,���\���[�Z��٩9�-�&`���8�N�G$$	q�H��Ɩ�е��"�`�4�Ul*�)�4Vw>J�e�Q9*�J��"��ю�V��W�5��G���ː �-T'򮪱�{�8*} 颤�/ۯH�:�W��9~��hG^3z��Бƌ����,3�b�mZ�7k�A?��d�TI�=�.8���v�����Wx�.�|K֐1�U��l,灴�m�{�n�n�o�P�t\�����fA�^� B�����p�	�H��z�7-٣����D�lF����w碤F�+Ky�6�f� z�Hp\�N��#0���͌�*3�GҊ�R@��rx��J�g��<S��}K�@?�si�O�d��'����#j��.�C��#�'`�$�[%O��e���;�������I%(.�T�V���*����xqa�>Ο�� c��w�����]L�*�� 6qL���x��d�i놏d�i0�^�L4���D]��ָ6M����)λdP���c�8��$k��$��H�%O��氻��<	��kxRp���
�V��%\_�Kf�0�A7$F!b��Y�G��¯E�r��	�ų
�+d^+�nI����p-�9�)�Ռ�́#7~��by	��ݺ�Ȋ�P,�!�&�D
�/Q�i��U�m#���Iu�������'���^EPN��X�2
3t-O�8v�L�qS��􊇔켶넏�1'$��'�R��K<#�d�����t�XP��+ҿ��f^1�Hu8Vݤ(���ېX�\x_��d�B�ʉ8-B��	��&Y3���X�J�?�Λ��v�瀚��(��K��?f�eMJֵ�/�Z�[��k��r�#����T$�d��ۃ(�N�h�R��\��S�Z���'�";�켏��э���������`��P��9�.��n�8���t㥅d�D�t�ͽpe�6W���җ��'F3�7�|�ވ�J����_;`0��A��4t�5v��J�@eK�o���N~�/vve�á����f�⳨�͡�vV��Qh9��_Cɂ�	I#;`-����ح��Ez��5]Z�1�{ ��-:P��z��4ψz�(�r�����F�:��23���n�d|�^4�Naچ,�P����3f�.5����*�1B�O<�0��H�Ff������,�K^��i5�C7�<�pJ�!rQ�i�+]����z鿱Ą���w�,��˪bm�e�w�܅Y�`�0{?�M�H4����� �S�Z��f��(���߻�Ƀ����ʛθ�iچ9��ﵝ:���3��9>��H?ÿ ���ɄR�4U�ƝC<x��O�A�NN�Ă���{�g�<���>`J�\Z���׬z9��n!�G�
HDȤ�����r
��eN�_��p�ӫ@E�ϝ��(�i�ӬU�D�gevgvƙ�JgC�ME0,4�av%�?��I=T�AN�8�2O��:�R9�#�~�p��SԠu���lP����~ݒ�'L�@��E��牬�vYK��nJj�;�*'�ns�!'�ѲƜ�A���`�d��ӱ�d��tcȎ����ں�iI�l�,���� ��\�5<p�cW�KZ�8Q9e(�H;�V�p�M��VY]��G%���q���\A
g�� tc �ǜ��}���<Ε��b}e!�T��u�/�;a�ejЗH�eV�N1r?�WH┥ì����䏝|���1w�\A��^��­�@�+[L������ �7�,'��ȓ��pU0/-IggttG���J�iW�l�B�7�iKi mK��'����J�7,�d��7 /,�Eƅl�M���1��-S\,�e�t_h4�Ú=�4�m1��NvbI��&�ٺ~�Z�܆\�7��t�SX<�ĸ���	åtso��fs���
�Ә��ͧ���ܱL��i���L�J7&�z/JRW��Q4�B9�'w��?��%5n��A������ڠ]9�`���iH s���A��	�Ơ`���E���.Y�ȼaL����/%��X��{0�`sPd��-E(
�)�W�*p V�y����� �f	�l�r�T�$^Ijܒ�v� pΗ\�$f֗�I�3;8��-c����c���h"H%����׹{��)8<�4�"��w͢Gm:���w)3Df_5�h!�l�j�V_Aw<����Y^c�b<�����h�#\�D\��D��H- �[�ؽq��ġ�Sg/���S�Z���o�;M��� Ԧ�-]���R��8^�+�$����f��XB�R$�a��$-\�����Bz���i.��u;^��;�׾e^E���y��y��`�h�Z����dR�^�飽�d�fh�|�O��vĉ#�,'J����������"��������6W�V�=��do�u�eh�TgF	!�p����zM��eH�ňȭ���[�o�t��Y����C ����#��R�<����1*e�[	0�A�ay���R{"ĩ�`�
?SX>�x�G�`�E��$j���g�`�����1���߽��R�� �d�T�)ǁ�=fga����ا�G}�4^k� ���C�'���ʗ(�~@\��u��(��Jˊ��_�Ӏ�s|�?"9���Z�F>���LBZ�U��DE���׊:��������S~��vK��A�.E��]+�#����a��O�}�)�X���T/�u6����a��X}��Z��]c�r{ކʋ/]�
�E��-ek��5��i��� 9Ǻ�y��3�f��ᙸ
~��_9l�Z�q'en���,�H�������-���6�2jA�!P��C��P鹐�}9Z*s��0,��I�����e�G�m��q�)��-Ե�\BYd}AnXo�^n�y'��j�Z}*dc�A�q�$CX_�B����{��٧���t�kO�j�L( �)��"�ɪ$bsR��'cq�k+T��R=l����}v^��>���hps���;Ëms+�"p@��,Kz -y�`����W���?�sG�����,cL������k�a�p��ixO���%B�!�+{�����h f�^�V��������VgJ������EN�Zj�KS�L��`��u���o$�qHo&1w������}�Ʊ�� nuT�Y<�w�M��P�W��t[����LBP��%�ٲ[DiIn"���熆�mj�a����G��/?�rQ�Ķ�s���6�����Zf���}U�hM;�G�?Ǌj�h[��Jȑ��r%��қX�r�y�=H��M?+�`�����Cf}ۭ���Z�l��u��)��\�����N�,���C�A��g���7�QƦm��s�*�~�ٹk���XxǗ�j�j�₨WjvW*܎��N%_���k�v���Sژ��u-Cz��^ٕ�&	(�a�3i���K�F~�:�����J%�".;�!Msi^l���?&��V��m�JRI���t��.M�K�E �z��ֆO�����7'W�Q�J���V���l1j;��瀎��qm�v�Ӈ����7G<��V��&��֭Su�&�t!h��=&oȢ��\������F����E�@l2�6L����+�e��]*	5S|fm�1�Ԯ�i$�*e�BR��,K�n�����K�g����`���ipk&��m����W�D��mU�uՐ*>�P��}�o.�7�%�)oǿ��`� �&��Xz��{�i����m�4 ��.d���::*
�u�M_���2˞L�#�IU��c�L�I����A��p��UZ��҅o! GS�F���ۆ�����F�M�@tGNF���>���3��8����/N_c���M�i��sSiB0 Ɲ�i��3�,W)��#U~@����w�-�w+��L����^g@���p���њ@�暙llH4�i�V�o�#ld�^2��8vUL���X�S%�f8�IZdH����)`��P�̧4%�
���v�e#2��ۂ�C?Y�q87�����a)3շ�
y-�������f��jJcN!Z��tȿ��6��3��=���<�G$�+�m����7��<�ۓ�h����oϔ�nU����x���#e�B�G8���G�CY����r��m����E���Ӝ�!d�V�s�1�a�YX!K�$1�֍Ԍe������=��,6:�qZ���9kSj,�;��~h�ݚ坵ط�Q�^jӈ�G�l_&��Z����wu�0�����T:L�1ѿ�?����k�S8��8�^��W��K�7�N;�vZ�(� ��N N�,ő]uן�b�����K�����L���whU���Й>��4����d��8�HY��6r��`P��S� ��\h�n����@d�h�1�P�W v^�q�2;D�П5qߎ�IK��$c_E�9g�[`�>V�i�i�Z�u��X�d���p۪�H�E�J��QL�>��Y��MkS�d
�64�vBo��C��Y�2����2��߸�$Z������mj9��Ac4<���N���[:���ɪ�}�ɔ;	�Z��X����!�a�Tr$��G��5�|�h��%I��&t�KRq��I�����}�(�Wo���30i�N�o���L��h!z�p�������J0����/������%ؠ��A����t|��h��0�ḲܐK]�.�s9�2��Gw�F��������L���dB
�P���:�f�2���b麌����{Pa
��ۨ'?�M�i'�KB�QT���@�9��w6����G�C��	b��1O.:�L�B폚��ە����ag�ѣrH+�����D��2ƴ�?���W��7ú�aB�	љp���m�O�-A��Y��D���:��Z��@l�U�7X�ӟ���w�P�����k���f�7�N�\�ӕ�]��j�9���q����N\M��,w�!��W�����H^�|�e^��}q���DQa��D�4H�o)P�~���e`�?uz���b�q<;��i��P	��PG�O~�.�y4wHb ��@v�s��:�	"��/��Nx�X�@����N����9�Vh�#�?x`k᾽�rk0�����R_.p|yI�$����R:��	Py��C*�u4�;�|'w��{&~ŷ�y�GK����"otc��/����X����u�+m�q	�׀�	1U�W��u�9�j�2�@���|��9<��R����ˁnp�5'�lpD4���E���l�\w��oa�Fv(\Dx,�0-�m���i��!�� A@e�e�a8�~�����[�t��ܥ/w�;���P;���ސ�����B>��1]���@|�6���Zo\�4�����n���!�~{}L�Q|��Ԗ�(t�a�A���58�3�967�!���R�l�N���W��R��d�hh�/zCU��2p��_���f���+�b�|� �?CA���N\Eŭ�uX���/��1�H�Ž�uP�_�z$Zxc�� �ppؓbP]/�YVP�������sk���`�t~ߧ��g<�wJ%�q��=�Ċ"�L��kV�+��nw������
U�H�䏘�2���
z�u�sÍv(3~��؅@����ޛ��@RIA������Z���k�.H�o���e��	YO�p�#�4�#��f݃ۄK&��q^��Q�C�	�ܞ�{�J],X���W��ĉ!�Y��Z�T� ��Th��KlDD�=ju���jo�vl*-(��s����C�L� �3U7���_{2�ݗ1�%��"�q�;�zd �c����Ό��o�����#ս�kHh�t,ZeTgL}��h=��S^�����I�YR���/���D�A"���k��t ���xC�X�{�������,�,�UY��$O����6HN��N���-�E�ㆭ5*�=_G���`Ӣ@�_sϠ���E���9~C��7�ɦ8�81�7zL��LJ���0)u�� �C���q�jӏ��<��qxA�,�K�Z�"�;$��]��a�qCw��ܯV`t��ˌ����O\tV��,����)7�`pbSĶ�uy�]��dfer��c� �[�As�elIG;�tr�=	R'`P��Z�"��Z�}�U:�=�k��\R�y��E�c����ϟ2�˾=M�xc�%�p�b�<ּ�I60=JI&��͟2��o����L��f��r6[O肰�r�+�kGi�	H�rٕ�HDyo;*A�a-�FfS^m����S�DH����;L������H��VM�ɀ�u	�"��������^xM���}��M@�DÒ{�<ʎ@/�[k�JN3o:\]�W�=[��k��gJ<#ھi�~>Մ^��JBp�w�琯�#��q�	��
W�G��YRr>
�͆;S,�fzXsӽ� ���WL���)�*t�$A���UN�d���(�װmq�$+��8n|;���u&���3��O�Ἁ'ִ�������@ϝ	�B��J$}�Q�e�̈�ag��DZ��T�����=Qc�����x��D��6q�l�*~3|�ƙ.�Ǆ�HZy�
Ω[�*�w�#��U�HySlvV�f\�ճ��nCt�a���3�������Y�0�ƉQ���7�t>���vFE�3���5��p����o�bA�J'���F��}L�/4s�̍�����%i��S6�b�8ZF�o5�1�6ق�Ӥ��a Zm�f�O�\td�i	�v��Z�?�ܷ��e	�qvXְ����)�-q�f\�g_wI%���\����&��1?�OGzb戧�@a�*��`�#ΰ���>Rŀ����Q����b�)�ؕ�A)h|X۷��5	h+�[ߺ��~��/�g��.� J�W�M�r�Qp�0���)Hİ[���x��adF�z����~�s{Pw�M�H���>�X��R��1�B+�m�âf��p��t���T@T^z�yY@L��F�)�����Zগ��
�J02��p?�캖޼�x����Z��M)�$�큝�+�̨���\�e�<R=���W��J�|9�f,;�4��.�O.ͷ+L6=f[��F�#9�4�f�|�T]љ0����x&Pt�S�C�`�V��ReW��CM�R��8�@��9ؾ�p��^�̃|�t�D|]�i�:[@����r끚�]C4�<���sޭ8V�\���u���>�替 |�
��M7��}��H��¾4�Q`� R'�>�����<B�/an��_ʱ�'�%�����
�!wp�������I�,�ޫHu�Z&���i]����̪���d � ��bE�4���= %��T8�3/���Z4C륾
��q�J�ه���6r�݈Kp';Lk�^Ӣ��Luv I���S�K����h�l:i�r`6���(X�m�� �#��Ig}�1�MeH���'8���qvE��*gG�Gkz�&��]L����ttor��!R'�aAʹdOh�Ll�S��>��]i�^`��}'��\�;�&=���}�7NC�W��Zh�J���P*yP��:������R�td��L��ahسg 0Aq�5Z�[Ѳl,��ύ^408!P"�����3̐0H![)}?�if�迲x��znC�e2$�r�_5'L����z7\�w{�̘`�uv�hAΓ��ړ8��4*y��Ϟ���j�u�s�1�Im��*��K���a�Ϋ��8і�|�y�_�6G4|5��V�,�dc��r��x�'�]�ޅ�a!��e��kn:�JT8~�	
��;v*ҙk����3��_�y� ��x+(/?E��K��%'��L<��Q�Z� ���6���VQ�w4��ڽ��J���������/���z���8���O�����^���P�X��V �Ď�5����~G���V'b}zZ!��,���9�,���i0��uA��0!��ѥ��$�4�S��e��ly$�-@W/ ^:���?�
;c��I�b�ߝ���������蔳B9�����++A��7¸#�Z�]G�G���&��z������=	2�%q%��<��s���H��������l���	�O?�KOR�42I�b`	l�=Yg��;rGB�:������q�����o0���CrOG�>F^���Ѹ�q���3�ng� �Hݼ�6']�}~���w�0��4
��{�׸�S���U�q���B&'m�b�q�<'���Ta}1NX�BeZ̛^z�7�>ۊ{J�!��a)1i\�����������l�Xw��~�ҡ ��\n���'f
�h%�ܹ��B� �E��+'u���P�v3og��$ť��������r��hS��9v3��@;r!�(P�{;��eho7��o��F���ȥ�u�|�+��|eF������h@G�9���K�
��V��$��u���,ai���3�ʗG�JVU����`��/��w.�
�_��Qk������^��L�]|.��I6�~EC�b��������~8�te���皹��=G����/g3?�&��~kgɴL�-���e���*_W~0�t��IR?( ^�PrqxP���������x%���L���H@#K������l��5��� �R���:�eTX�Z3�4��a7a��Z.��n4&�@͟LwQ�71[<��~c�ft�M�����n���%&��|��^��m����Lݖ#��g(d��+��g��<?�	�АjB��*ǋ��}��\
�tMUb�!n�M���W�i����TZ�i�t1#����َV�M��)��K���d�L���i�s�ēԴJ�3���"eG������&��?�{��S��*���AX�.Z�a;^�e�[IK/�h����3  2���+�P�d�=>(e6�O��;�o;�W��}Ŏi,��d��u���M9ȧ,�so��s�N�� ��W��wHu��ͪ>���y'��̑���\̈|2�>l翞�@k��K�m�ȵ�_4h�����N��!���R�ӫ��ΌJ��x���5�ߛp��B
��;�8 �U;�ڥ�M��讆�\T����(O�������}BEJ�2��sS�x���|V���Mu�/+,�8^�#��Ph���J��ИC��8\�!�IY������g��_s�'�53����<�{�L��Z׉m�����u��S���M&;h���S�'ȳ&�Ip?-+75L1Hv�j�2�!��ۆt�D��G�� Ҡa�X?�ۓ�ehrr	���E�v����6|Hj���q?�_����K�
�M��N뽬�S��x�0F���y�����D�&3��*o�4	/�Uj|R�G���Lr0��=^l� �X���TxJ9-�
R�o�Q�	R���<R.+��~&k��J]�T���y��`��H[u,UQ���;���a�8���U��o?�c~ nKT�Hx�8��d��A@
"ok�Ij`!��s���(��Ay���������bc;n�N�'����� RB��0�H�<���lN�X����?8;��# �:�|)��$^�r���#�}��E	\�
G����6Y5V�C��bn+}���F�'ĊC��e��r���W��vS����d���Y���,�q&b&N�4�Bq�����U�M����I�@/�rr�ƌ�$�A-�����z�Gx�����P��J���1_)X #K��@%��m�YN\� {W��WP�F���d:��E˻v�1#"��a�H2-A��KvY���6��S^�`�-��,�L���)�1 >�󟤎�m���(	&����F�a;WHN'<��Ĺ��mIS��X8!@��rv��l�0w�9��/���Wn�F_SAh\m����AҢ��p�ҝ�k	C�W�͘6��d���㽗o5�v��4�@���nZoV�M�8�Z��;�h�V�IՃ(�Ђ��:k!�d��F,����V7z�G�O}�=	��V[9n���Mc�H��_Ȕ%MǤr&|OS�]��Vτ�>���F�'G|����U��T�-i�����4$t�2��I3�:���zDP��R�/S,����D��A3~��|W*j���ֈad����}�����x���ќF3��!�B�C���G?�rT�\���k!ă`��� y;@���d8�y��o��(Yj7�: ba�5�U"iל>��
k �S,�	ӱH<а��z�eւ͚�j�y~����&!��؇oϢ|>v3����z��j�e��*W)��3'��ʹ7�?��q@�[�D̓���i�K(�����#$q�������r����k��O:(��;�V�j���7z�P�LJ좔�G.1w���t���҈�ӟK��������"oo����4��Ϋ}P0
,>3�:rFǕ."�A�#�wHz� �V�/h��W-�>[���W.��\l���5���D��60���T��щQ,u��N��6����+�74N2�Z�)VJ*�d2��ĴaDi���":�.��Ў8��Y��\��S����efnC��C�"*��#t�8��v*�Ns�Ca�	AM�q(C����ȴ��'�F�F"�#��W%o�H�PiC�6���J�D�ۤ�S��-1\�@�߾���ѻ���\���lQKv����
<�/�|�uO�Bd"�Ն�H�f�\$�q.�ݴ{������%�ɍ�����	`=��\CQV2
Rn�݃~���Hi��y~���ϖf栬z#5h��į]P�_|ܑ^�D-9w����p��>���~��V��̷NaK�EWv�H�Y��!v4ô���}�"���e�V�.4cע�ã��x�^:����*��>c����k��.IZh���7�emH���\�;�\0�xn��I�=ZB�xNd�Z��a;��]L�8�ƺٚ�u�%'UĞ��Jan��h�o�l~Yt�J��?%�����/�Zt�G] �H��k�z��j��y~�=H\4FD�K-K�h }�� N��G�"h���|���j%ڰ�84}��u<tX�il)=+M�m
|ݘ ���e)�c���dKO�|>5<_�j���q{�iQ��v1LҡF�s˄�ve�O��UV6��\NU�4~�_���B����
�-��K���`����bx@Vr]l�������*��_u0M��~4<�(��i��M���b���������8#9�%c'��ÿ���� ����jIT��I���r�c!f��ҋ%���g�u��E޵�sA2�F乡�7(��?=������|�_�{,�"oȷ� �:s�r��L�M/~#G�|)�����ƙ(�is���
�-���(g\Aq��iF�QOV�%�zh[8賂cO��P�Q��L��$k ���k�]�nd�F�v.Oy�ll}��Af�����6���o�O�9�-b��v�>����tm�N��ݙ����p�n`_��E�z^^��?���C��g0����4䉉����	rc'��f!yJj���i76�wj`3rƽt���;�p��@�!�Ty+*���������I�EWj�`0��D�_{cr��Ǒ	n�}��9���?��Dh��b�����K��" 
�vH+��K���ho?T<�NyV��>�+Z@?�;���T�)�^��$X,�ޡ�!�aQ)��g#@��V# �~,�[�.e�tޥ�;K���KL�v<���ӯ���%�ry�����@��oY� ����@<K�֏�l�)�Ԧ�쾱��&�-���KJ���T���ɒ�����6�%Q{5�d�g~ڐ���:�q��P���63j?-�xX����fk.z[����/[_�c�I�;Ŗ�}r 4C��r���{r^/�m�h�;��!�$[b\���zV�ˮ��������ʾJ;�I��\fY
a}����@�[��,%R�h��p#'~w�<;���a�2�~���1`��]�T>�	��ۛ���.&B����5��k��:��)�L?P.�ѻͷ�i�HP��W��x�`i���HN~��L�� l6z�#9���t���e��u���[m-[����P����M&�A������HC}�������|���E/�9�G_�Ex�f��d��d�zMf���K���P�~��Y�^�c��К$���9\�Θ@;P�40�7����CJ�_-��w�[ �Њ �ڬ)��mێ���XG�����_x�~�K��|�)&�Ğz
#�Xj]�ʫ(�t��d���YZ��ŏ�@v����� 	 {��V�&�J�?�	�kV�#N�s�}-�����������R��<ڐP���]��IXByh#~��B�(��������p�������`=���yQ�JԲ��SQ��>��}�,�z*�:���g��q!0d
�c��q��}E�"�b҇�'�x-����E�B�GO��^PE�<��㏽�!A��O	xr]J�	���lg���N���Ŀ�7XE��)�|��A=a��6S����&ׯőj@7�\�����mJ1Rd�������9Ll���� }`%�kS'�P��-+����gnP��>���V��lurryn�������+��A���[uN�Xä゜Ow���MRz|A�lȼL�$�`f=�ӈ�����,�{����g'�>�z����ג��]e^��h��:W	�<_�B*��<K���X<v9���L:۱f�Н�j�����}0O $7�M���֥r�`�	~�MF���%Ǉ����=����5Ld��DzlN�v���3��K��IDj�ҁ�0AT:�g�E��1X�"��<�k���.*˭�����k%���˽ȯ@Ĉ"B�0��F�U��i�%�^�������A�=�=��K$�n�����(�Q)9�v���]��.�"4}v�[��ow
`B,Q�|;�����fH
��3j8WZ���B�^%�ʶ�?�UX��W ��Cе�v�%�����rY�"-��],e�������a5�\�t��`���[�Q"I!JE�$|��l�`���BX�b�,a��W�Ax�Jk�
U���o��>�`���h5�S����4R�0�b��8��Rx�y���X�}�_�������O�Re��ΫY�K%q��[���_���4��C��Of]� "�(��`o�2��5��F47�����9��k���nt���2(#��i�Vu,I>4x�22LB �v�P����pɬ�s�=NW��7�VPfM�6B�WZr�N�p�۾���D�4<�;EyBM5�d�"���XF��!5\���u�a[y�����@�fT�m1@k�(�N�%.��c���#��I�m=�{�ՐD.��j�3�����GY�ua���ĝ!�\[Z�@���W���o8����c?���%�Yѭ�|\�������p���௯����P���(	d1�|�??w4�r���߶^��e�G^��d�t�!��b_{N�!�W1���6��.�:���=��E$j�q�w�r\��r����M�������nnb����ސ�����[���${J��cW��˟���F�)!��Ky�2�\qx���$>T`��j\���QE�`�\�%��c�^�ϧ����lc�(�G��É�-^��5�̴�N���%A�<تe=C�X����r*Y�ýM��#9BS�*5��C�C��M���\>��FGƬ9��v�ʵ�M�Ϙ7�\W�� ��c���G׷��{^<�e]y(>a~��e����T�H���ĊQ7��Ŷ�'/Ws�Y�n7Q���T�FXs���,�LPJ��.��� 9A�C���'o�yɢ ���
nȽ����­Q�����`n�Yv�p9�}dH��C�#�ɕ݄�I�~����tS�����@<��l.�.����r�°#���I�N�A�u.v3\���V$��+��qD]ۖ�t!P\R��s-& �}Y���/2I\����"CJ~���-��$�])e���U��пd%��_��Fٚe��:�:�FQݗ�; �7�[|+�(2}���<�	��),�׿�_ �#�yu\����Yw�}�շ8�J���!���Ede�J.���H@AK,Τ������<�_���pcB��_t`��>�^����g�֐����լM���5�j��O���?��A�}:���/3j�mG׹�s0oс�r�>A$(u4T��L��)2���T]�4�ػvf+y��L3ތ��ߴ�&L��[*Ճ����o�K�b.���}t���r���_�΁�=Gu�^�o�����'a f�Τ�v���.���Y�l��ߗo,��i5ov���>&9���[~W�$�w�Zn#���G��?���ʛ�'�]y��jq+ש?�;�fタNl�i���!�ĝ������Y�1���T���l��A	h����wWfT��N}or��ybU�ߐS(��ùڋB�DC��2��֌�Қ�)�Q!}�?�_d��dg�����[M0e��*�O��-���@-:=�ۨ���[��V},����<h�.YUv�[�2<�9�"1�wꜳ�t\�4\ӀM5U��t�2�S��wG�|;30ʬ�r�����0%�7%Ym�TvY![��5Y����s��x)�z��df�õ wd�Թ r��.�P���c�%֬�{#xf�hb��4���*�x����0h�*06�`I��l\�kR:�:�L��r�7h؝Ǥ)�^���_�n��S�Ӆ8���	�^zv �o~EzYX��i"Y�ר�h���f�A \.�.��"}?��`�����Cog"��[�>�Q��։u�'�@|Ď���ԃ���Xs��>��=�q�X q��
Ə�N'ȳ2O�Sa�u�����q:�s�u���§��쨩o����Dm���֛3|�ʷ)���g{E�o=���F�M�2�={g`�r�7�]�~N)���d�xuFyJ!��:�B=va"H�h��:1\쎺)��;���ܳ�d�h���_���1W���|$w���%�y7�=Vd j�D
>�5�~����F�^n ��F�Dv.(��cAƼ��"*��G
Ҿ�=��6 ��X��Z��V�	�ڙ���y�:c�6@</Z�Q�_nA3�	茨5�26�^��"7� �O�B��oG�!m�گխ�y�G���h�*��|l~�:5)��
���w�	���eA:�W�'�KfG�k�<MO��w!�VL�u���	1���v�nw)��{ެD���I�ٯ���ǃf#�) ��*'p`����]�<4/Ec7!��bתxJMp��5lؚ/6\�PZ��u_�$a>N-�w|Y�U���z��B�	X����!��D�i�7iz.Y / ��$�Y#���su1w7`���l��ۊ�,������s�/�����Gs�{ǁ�I��dS�d��	?\x��P�0FZ�98bFC�}�K�P$�{�8��i�?	S%������RLn
rY}]$�,d�o���-�Xpr[z�}j1���M6�����N��`�����['��g��8���[��Z ����V�O2�}�k��	���&��*x���{��奸�#�T�饒#hW�폯�����f'���P""� ����z������3_zn!O]��ɸ Rt�F����]��M�É���)��k͓O����j�)����$��|h�rª�,��ge�:��0T�*��S���_#5l:^����N]V~cD͟��������%V�����Sָ�.(���		Y���j]��5���㕠ZYl�Ņ1ę�WC�I���vO��~
��2��|u=�RV���/�`J���
�_�tZ@��+�ҋ�Z�&;g��lWD�n�J[L����O��nN��G�h���!*�\�-����������y�����qB�����}�Gg9y�L����3G@��@���\J&Jo��������5�_����v�񥛝�8Tikl7O0�����=v/��;�9էޥ���ՙS��G�2�+��C���Y��	����h_�H��V^��18�j���!��!P#�����J���P�9=8���J
�i�/'����z�aY�5]��)���G ��1�>8d�c��:�dڇ9*S�L���6�m �:;�������>��h7DR�֔�gA�����pǺ5ԧl5S\n����k�a��%�Df{�c�C�ToC�NB�6)���|D�+t6N�9'F}K�i�}�'���@�6�?���1�֑�W 72 �	4ʱ[�w�>��(4]���w�b��b����:o-���*-�ͳ��f�J����ok�I_�$�~�dљ��!��^�e[��wuq=*�'�*u�`�+k�tln�32�F�d5��Ir4܀O�@�/����uf�ށH�c��i�q�u�B}c�:��X��]M��`��6̀�T;�Qo��m�I�@D�Td^L�ze��
��̌v�%� h�u$W��U��Ǥ\��}��껣rP�٪��@Ule��ӔV�Dތ�����B[�a&R���^8�͗���W0�uk�^r�T%��43c���/6̖cv7�>�/�x?��R�l�@��-M�v�3ؠA㤏h��<����-��QE�;�0hXXdˬ����)1^h� �A�j��4�C���4���~����&�X��4�4꘶Z�GJ���+(a���;}�t�Q�&q��m���`���Ad[~j[>=��E9Z��ǓPi���;��m|�ڀ1>޿��*�N&sB���ћ����$�|�$i�K�mG��ٟ�����1�#U�b�X
����_�����?},��w��酬���b׍�!��w ��7=eF=f��I4�Ѝ�Ő��w��$7���@�$^��j��E�p¡�E��x�{��	���K�= ���D�@�"�d޷
��'�F�%�F��k�U���*��6� �^ �ό��e��q6��9Ї_�{ނ�ԃڣ�q8*!F)$T"B+pD����0)i�v&�Ր4%��������J�#+߆$[��)�����^�Ϋ��U�U��Z��ވt�M��kys`�g�n^yñ��l��Cnɝ!J<hJ5���ik6O2��$�:f�ܷ��쾟�v�Vq%�Dư4�"��m!�s��1�'��K!�xpB���uHm\Y�H�qFGB���ʄ�)�gFh��|��쫽O�J�N[[�WsI�>P�>�r�mj�"��Zy�~�j���O���8+|�[��׵找��.a*8�oIO���i�+�-8��k��O1�:f/e��1�	#oY�;�U
(�ڊ�{|Ss�+����x)&�����������ӷ�[����� ����T.�\��i�ć�c�-Aü@ �w��3T?�r�� ��JS���t��VH�X�uaٜ�����m���!'7��J��e���)�B�&# Q5G�t�Cң����"�oKN�(�?�i��HpX�lbo���'���Sn3�K��6��Ozi�f�EnD��k�ֽ�O�ti,2a��!��WA�S�{���R�g�"���/��VP������Ry���Ҍ[���Zf�N��d-	�N0��Χ�d��W�V?�!�Mܘ������ץe�+B+c�(����H~��+���ť�)���T��!�1�~�M���%[,�0,	�O;@��i��-�W|��brg9��c5�^~�}ېo��=�E��L�fa8�Q������Gezf�W�?	������X�4���#��ڀ���"Gğ�ͻN���k���F��.s�J��VL#c�2G�`�H'7ec�{9��~5�t�|)�G����s�ֱ�/m�R�K���В���lD�mкZP� �ECQ�o�ܙ9���� r�g%�ͦǞ���iw3����:���8D���e�� �h��
��kE�j8{&m�2�bik�����%�t���x������KMJÐ��4�K��n<�����f<Č�����E��Zp��;'g��ުB�$��<D#�K]ԩ�%��,�� �v�����ܐ�X���G��������'Qڀ�1 ßТ�g�f;=kzʡN}�����(3-Q�W�z��O�?~%?	do��BCz͊�|�#�e89u�/� ��6��;^![=�z�2 �?�Hx|·s��T��s���1�e.�wH�M�����_ɖ<�1�Gl��PL��[:��U�%L%���=��O��{/��q�9�,k�����g�t�t�� ��Ll@Sy4&�˟�#�:jT���D���{C˜�}Z.z"BQ��X��H���}:��;��|4*����"����v,���,%D_S�U�a�Mf�<�t�,�L6��Mg�;3!ˊw�L0l��<S26��1�L���V�2rg��;�q����;0 �>���>��j;��b�*
��qN�8��G=��W��B�q{dnEh<��ȁ� �L�PK��ts%���l7�p,�	x��)��b�R��S�|}}��{�.Z�AH7O�|]���9�A��7K�����H+ ��ʂ(�5�Ŭ�>��%�X8���P��P5�M���LK��< V^�u��3��u^�X5a���g�<�VyU!���7~����-R���ɍS���ۼ�ZA*�o��O%>	�g����0[ �]h4�3���Xz�p�sh&��mb#	��U�}&;|�Q�����(���� ����уA���>�D��x@�b�_�j4-�
S��8%}��Ga�G�ҕ���QH��}N�g��i�NNs����޻i�2�Sl�ɜ�7].�Z-��;O6�D���&@9Y߹�������zO�ꡲ�£�&8�hFm��#}'��N����v��ux�:P���n	σ�'�˖��.��n%����\8j�,�P�����w��,��I�����\��h+��h�dNg���&�y�)] �j6�on�{5�m`c���O{����'���'��Z򭨬p��")�BޥMjs���?c ��F�͊�N�"�!��� k\�q�O��s�<������6X���8.�+o�,	�:
�1_�xD���D}�f����f�k�j�$LP,�`�%��	�鱰��i�TO,������J	ܬ-9H�GE�DI��n0�ߐ>�����'�eA������{��tW���Gg=k�ˮ]UycdK�o������W�B��tC�BIB%>F×��B����:�k ��CU��f)
ق1��,m�[+xJ���}���(a��Hg�5\8�\��1M�o���	����w�N�fuW6�x`2~��0|[$U���	<mp|ҟÜK=���j�����*�z�3a���T����ƣ���F��܍d��6>USVy!�+	�8�RO	���hE�3#`~��x��3����&T�
줣@��J��B�	��hZ�}�zd[�n����v�1I�&�e�7���v�z_T��C���K!��M���pޤ�U�F}��!����.�����H�!d�=N��2��ǆ��3�sў�7�,PEڟ+��*QS�0N�$>>�
�'��1'_�$o��{B���|��s@G�F� �~�r96��P������؊]��
:d~=�x vu14�(�5��XѴ�;J�baI��8KO��+t�X^M	9�1i�g��U��Tf�u�n?���`�3vn��$F����jm�F�G�kzY�@
�m�rv�@�V� r�i㲰�9��@B��Wf�T4���/��D˶h�R�΀�TG���9��q��?LtO/�^���56�I�1�����J�Z��ݠ���h���m+x�)d���ŉ�w^oH#�$G59���U����L$l�n�D}tJ�$���4�y�!��0���::~J�a*�=��=S?K�92`F���G��ݿ%_<�7VJ���^�
f�h��+���e0���:�r��5��lL�c9U��ac�<��+��� �' 9��N����M���@��׺�n8����ޘsik��a�0������Z���^6F6��C!�� dJ+��{w�&���ʹ�XN|��R����2��i֮<�w�O���(��ydF��	cH����"ovi�@���fIK,݂x+�kvLz�w�{��[�"�m>6k��#Ab	Y�d%�LfT�1�/ƶ�h| ��R�U��$�g��0�Ak�M��˱�|����Q3|P�u4�`�������Z$�������u M6%Ѱ�/'��|�}۾��'�����B����@�u"Xgw��	�x�	`g��:��&̔�u�EUFJS��l��%����0�0�k��u�옏M�pQp��+�,�r<6�~ہ3O �Š�F��Ӯ�8��G�
B�K�"T�+ �O�Nt�,|@?���{苟�[t�����AёEZn�%�k������)p!w�6�%Yo&���0��������)f���0S���Yqɡ��//0�V�m.�u�'S�M����\a���k����Sf�Ԃ_�ڜ:�v�p�?�~F�ƀ��f����s�^#�_e��Ǵ�n'?���2P���ـ����k�iyL����&u�!m`�i!v���� V��Z_�P�!e�tCZ8Ҝ� ��_��j�� �wo�W�f��$J��>��K�a�d��H��5VD��R�q B��\(����XNJ8CLT�M��A��WKC㏠yF�'�;d���fd�뀀��;���J�j'�ap���$�Ņ�U������LK' ��QG����� ��*��B:I�Q2|��UUh��b�}�q9���Ҝ�Ђ�)�2�?��6qD�&��䴻) W$ļ���%��y���� �cq��Tz���	W*�h����(`��T�+\�V�n�n�\�:��4k�Tv��g{��p��,���~a;������+�^�w�Jz���_��u��8���Tˍa �ylH=ܮ�P���ԂVO~�r��P�r�ެtH�-�V&О�+
�B7=n_
�@6��d�0�����?�0������1�%��� ���e}���:^�ڬ�����3?U-6���<��M�l�Y�Y'�m"#�l�����pg�&6��j�w�*�p�1��u:Eh��/�r�'M:��&Ua(��)k��.���n��+��#�9�N��˲�Ꝅ^�_n'�r�ʊ�ET�k�t����(ls���~�`���{�}�Ej�"��1�^��ӽ�؁����@!�W�ղ$�v	�f���b-��:o�P�3ˈ�g1��+�j��0����h"(�e��q�����M��ѡ>���nk^�����"U#P�MKI��T�0Ҫ��	�E�o��|=�`���t��[��������z������ܺC �j�	WM6��N�5�v��(��p�y?��"QqH����29	��#��Š�����*f�c��Rʫ2���+FUD�d��D��IO�`�F>JZm�$�O�]�Ga�%��퇲�]��w0kKs�������C)C W�$C������e�˭�X_�/��Lp��!�Q�m9��څ�)x����Y���OT�o��:z+s��!]̺w{�NR^�bX����[�Z��-� �D6!u�zJXQ�*�vb+.���,��-K�!�k;"Թ" äwtow�� �_p��zlo�y�c�k]��`f�8�������r����Ow^���VXj�8C�R�O�Mlӎ�� ���<,���c����*Of�� ��@���_Ĵ��0�;�K�$��T7���,�����}+=�M#1��z�!gJ����_f���*\y<��K���E�\��fj�Kp��
�'%��W%�~��Z����L��"[�飝������r֌뚴�3�T��ozd�9o�rZ�����4�`���F�1:h����1L�E�dÆ�K&�-t�F<X$�y5���� =ɟ(�*/FDx�&�J/8�Bkuտ�����Z
��尋�����'�5/,��w�P�|��|]n�cE����W�!���sk=�WO�Ӻ�	��p����zwy�ٵ݇��e��Y�Qλ�E7�OheE����n#0��: �o�+�M���H�� �KR`hްKB�ky������艁��d�ԩ�;or,d��D��;_VF�C��5�R���Zjk��֓��"_Mu�@c�:�������`S]��^o]*?/W`�W�0��v��z�D��e �
���<XY\�<�k�n���	f��W']� 7:�v�4	�9�%��J� ��?�}�����M��{f�w#���V>�j%U5ޅ0>��Ȥ9^��H����7��`es �å�������Mz���!+�����I�2��h��}���0��b�v�v�x��Z��js�t����xP�\;�*z�:љ$!S>��c���o�V|�k�;����䉰�0s��͖M>��(pT�iնBJ�s0ٺ\�����Oз]e�x;��ոfo$ ��4���T���d]nMť�����8����`�d%�;�_����[����)�sڥܐ_�*T�_pX_���eP��̘�=���fo���ПC�e,��pV���������c���;�;[�bm�N&��׹.J���FbO�"z�G!��j�&0���Q#ƕ�K�Dw*���6��4�5�SX�h3k��1�'�ˌ����%fb��mH��.*��2O�+��6qv/���BN���,$���SM��LU!��� b��z}`��[>3C<�ZM[++V��XDBi\̡]���#�c ?����ȅS=VR���x�	c���X��{Z�#��W�d��em��ښ
�����i'~�ة��JMb�t�:�}��c�9j4SW A؛mǗ��)�V�6��
��|Cm��gK��|�&:�b��]aq�#t2�S��!j���݇wx�Ӣ��&��pTWy�`���2M�P]K6��L�����MzQ9�Zm]d�G���f�-�8���Ȼ�IB�{q�t\dFi�b���F�1�>����+r۹d�T"n'���Y!)���ڮ��\,�'�H�Ģ^P!袉���G.M*�8J?�@�� +P�p��^<{�o1+,�����O�,��R���	qqOb6�����"T�uQ�t�o�s�}�9۳�}|���
�'}�!���|�d�&�����#q�\�����d�������>��!�(Z�y���A��"��Xp�QDMP��ӭ� ]`�� � �������q��ZUR���Dm!4[�M
���ڄ�}Y�D����j���0d"'�ɒ���0�)N�8W ��h%T�ݴ	�zvƖ8 ��֎��e��Z��9]eE�|'v#i��O����O?z��^�S�K�{����ȭ�6F�]��bK5�8��`�Ou��:�S���D8������p8���$V��;V7*r��ҽ@[�]T70V��)��b���o	`j��?��.;���ur���ն'oAQ�	Y��g3�Ȗ[ur�m��p���/�������%�Iz�Q\(�Ō�#�9��m�w�o� 89x
1���Go%,VX{7�Z��!MD���%Z��zi��O������hdt�6�
�p��U��BcZC�Ŗ�*:� ������RbY�9�1:=s��Ķ�"�/W�F�s?%���!{��|a.���N(p�+��u�S;@� �����@��XV�R@<�Ύ.Z!s�s�3T�.?u�T%rg_��Vl6�3���C�a��D����S��]BPx�ea1I;M����Q4�Q�Ϟ�*��GD?}#[44�����*H��';�G%��%M��9�8�� q����fԯ���q(�k+v�۳̥[��y&z+�ۖG^}<� w7n���]�-�?s������*����e��3c+�Or7T'&���N�${������;�>�J�uѳ\��5�J+J'�޵�J� ر*~f�A�$��M4<��A�Z���Q��a�������;��UN�>���@���V+l)�v�R%a�)S/SVr=�H �U~쥚NJc͙��s/<�3�!�7Q����B*�p2�Y�W��Gc��ߛfʚ�K��Vq��&�*����]����7�ڠv�:�U��B:��(��o���<��{B��Ec%��prM�֔ީ���	��fw�j`�]��Ó�<2Hc��9��]�sf�Bk��������!U��2Eu�2�Gf��"d��YfbC�y����5���3����SzyY�W�6��[�6i'ɐR(�k��d�-�A;��W��6p�NS�M��'�Uԡ|��Bֺ�d��t�:֠���r]a�����c|4��V1W�%���E(֬��q�~.=�!��i�V�ג�8�\kܳ�s�n��~�4���v�va��^&Q �K�|cD�p��X���语i����u��&z�t�j@0�!���Y�m�����\1g��@�.�a���cCx��T-I��Z�ٶɖQ�J	���q^�������T��@�@9��*�e`Y���f>lg���n��>��'gH-��אY��ЕV�6�������>�j.��F�f,k�w��X�s�ܛ;��Vylˣ]��F{֧�}��)��ז��n��q���0����&7�La=�D[N�,���u� y�=ˮ�;M~�I󺏝��U�k�nH�R�9?B�
E�dE�ЙU��&- �W�&�|��F���<w�6�'��Wx]54_v>x��y_0$�mXݶN��zS���@��k�$V�����J1�����@_&���҄V����D	�XKѯ�t_����yI�7��`b�ja�Ӄ��g�X9���9�Ea�t�
��\"ʄ@�a�ǐa]���~���gf��þ�7���1N#���vP�Kd,�GZ��l�q���ۋ��D�B��j"u���Z�q�ȭ��p��d��<e˩�]�%��R�+o���R��j���N��\��Y�G����$D.���y�%�����h��O�����c�"Ch@.9���}D�	��*�VpAq��*&�^�i�m�$�,	�5�}�E3��(��䎷����MoUf���zՌp{�0������E�c�Ur��]�p[���u��	�D�c\���T�&9�[7�����M+�U�z�l|����V���Bk~Mrk�	��͞��r��O�ȃ�<X����NP�/�Tޞ�����k�WJ�h 2���m���fF�`�4�wG���ڹ=v���U�7�J_�t/��X7��F��(��R�!���T�;N�T*�:2�&]D�7���f��Xr����^*�1ȥ��Fx�?�v�x>Sf�Z<���*������>q�M\�Y���.Ce�
O�l���o�;�_y�r�d�v�r�?lBxՒr)�ն�.��������Qn}8�T�J�s��H&~6%۬���	�{M,�]V�=����ô�Γ�t��{K��Nd� ���AP[����;w[qx}�`��ݻ�=����Ƈ_�/���|�)�kF�������F�U]2XnZf�l���%}`c:��������Ŗ�� ��ڈ���i��.)%�٩�+eÁc&F��K�*&�����ܕe�{Fl3u��PC���N��9(<���O��oO�3Ġ���t]0:M��m��C�,m�͌�ù�8�����c�I���@{ӘJ&\����� �"��r�6q����	̘:�Ɔ?��Pg�g)��T2$�S� V, �c����]LD��;���������e�m)�[�x'ĢR8/޼!�9�Kv��3��B�9|'~E����B�W�1ծ�o�=�>}c�s�������yk5�_"��bi3JK:�wZKH��pS9�F�`"wz�c�"��򹭜9Sk��~�5���}�r�2dLm��%:���S@ӱ\�@�l���MY.���(���Ƴ�4�'ڏfa"��r 	�
�ƺe�笧���V�b��um�<�u�
�\_��zN�	�y0��`h*���kś����2{mQR����6��v�����~�nMs(\�9�lTs4�GE�[�fH�f�6����s�C%E�
S��9��\�po!C�rJڠ&f5FC:��b����� ��
���*�[S�HKg`%b�qY�t�V�����8��,�>]5\(&�)/�ޘ�4����͟/~c���W�*]*@5܅�%�j��ꈋx'�9)S�t�*n8C���Q�����ε�X��m���*��`8�׷L��CVe����m�^'��K$�3�[2����U̶]�_�7�F�.q_�'V#����;�&BO��&�f*��@Ֆ�N�/��je@G`$�P¹1�{���%ό�w�E�����^�}��9���:�ѹ���������3wA�~�'�^+$�C��� ˚�$6����ϥ��$#�1n���~�ȱ�H?! H�5�ܒO淼��v�%�o�V=�:�m $�5H�:����p`E�1Ag��i�<	m��k+��@��m���a�|�]�NOʃͲ*�����'v�kƬ~���@P�q�����Y��Ե9�P�W=�j�,��Xz���z�LjO�"�3fKAY����������,�ՎC�`��*c��7!�˜2d��-B�/#�v��I����%�zz���W(�x`��
����r�%}�����+bEՒ�A�� ��u�x2���,�HB�w�D�S�0��]�$w�:��ڦ�}�c �s��E.(��,Nhc��&m��EBQ��X"�'t���g�G���蔢�`�\�Oqs�:�뛷D�j�v�6���٥g�%b>�dn�<�%f���M\ڽ[-t��ן>�MQ�o
1o�l�Q��ȉEe�9n$�Y}L�����	���2�S:=�{&�y"qA,Ѵ�9(_0��������?;/v�U��#�d�l���): �g�x�u��x�dn����=1�
�:B����6��E'{�=�;X���k�B���F�^/�ig�íQ�7���WNֆ<(9��	�۫�;#��QC2gv&иb2���9'Q{|��F���Ϛ�+�6���.?H�T��_Ͽl0�#4�x�:�~�T��XJ&�=!�f3�Kb������vGf�������-9�m��^��ft�+ԄLJ+��ʷ=}�8ҷ�
_�b�.�ЃI:����Ou�
;3��C���6�.YG����Q���S�%H���ơ��?.�V����ֻCC<^��%�8��O�H��.�?�W�Ϭ�sg�<_�k#��,ƪ��o�K��
o��/i��Q��U�ZE��7,�%�5����9ef���ӠũV�^�:�@A�<hYh<�B���Ԡ�Ě05R���wi�L�*��uF{�I���y��'V�u*P�Nu�D��	��M ���A��q�4}���������1�J�&%C�M�6�?��_�$f���g�dg�|��ߥ��;j���*�1�V�6���f�T�tKݖ#ߗ��o1I�c��X�ӱ�T\ޭ?fd5M�[je��8$A��%?�l9��\�QH.��}��4(D�N�f&���5C�(��ZL��̥���\Ls�W��C�p�rv��x'����G�-"�l��kJC]!�Y2�ӍREse�\|��=���Zh������a6Cra��3�{`��veDwG>���h��Q{�M��Xg��n�4�ڽ��c������.�yK��>������p�#����4���.��"���h�僯�c@9J2d�=@�	�׋ԭ���c.���Fo��W�/8�������� P�K����Ĕ��`b3�ou���k�u [8��R_���G*�bz/���q�XOtH��W�/�䠌����&hGh=t�a��&_��-c�QRXq�~�[����.���'�=l���~Qsm	,��&��pI�9�e���N"��:.���式��m~-^[`�#��EF�#P�};��81��%�B�q��[F�^d.z[�]!P�pO�� �UB��Y�����<C%�􊙞r;��������K�5���T5 �UҾM=+�����O7�Q� �^6}ȴ6�����bM۩P.#X-f��p���u�*D�o.OP�&�=^9L�]�W݁�.��${Xwz��������ʜ
ȩ��w�ȇ����7��)/��ݣ~�BcMf���RC(Y*��'ݥ�Y�UX�i�8
����^p��q����R�V�����!�s@��6�nP%� `���Մ��s �(�6��/P�*� v6�'�J+�^-�V�S��2�I@��|����z�n��x+L�%��A�Z,n���x`�	�%"�9�O����2E.(�b�&����͠*�i�e7jq�27R�"�s��YQ�Q�Ւ���N�R7�X�_�
I��|ؓb���Q"��>����Y B�^��o��-��%�_�G��� ��q��X�"�{��ֶe0���Q'�-f=pM��b�<V���`�ck˺!��*�<"���qU�Nz?�h��%�G`��/R#��.��*#�����̧nEM�i�YTަ��c��$��5\�PB�\#t ���*�Ux�α�4]�2_2�R�h��WHAL�d���p㰐n��?[D�#�\�!Q7���I�����E���ۃ\m�5��#��"�l���Ь�m�a��d���[6lq���ǎ��}%h���Hf[�y��h
�����0���B� �t^���{'j5�����W�]
-3[4X'�P��uCҍ�M�;���r^Jkf>�S|�W�yK��&� ���Wxu��i�Ĳay�K��Ӻ �lP��*\��$j�_iH��J���L�^|�x3Kۢѩ>�S>(�:`8�(T`����E��Z��t
O�v�,Z#�4�3���Fi�E�P��f6�� �����FkK�1��%�k���i�>�v��S��n��3�z_W�N@!�Ç�K.�|d�+���H�1���W��!@�RL>�|�W>�sD���p��OC���@5ƚ	7P��'�����t��e,n��(�����!�kDGNLJ�x"t��Ai�2h+�0HU�Qv,�
j'�[�{�+��.����f��~IPё�'�����žb��k�%�|m͌@�,�i�V�f��1�I
6N�P�-��H��*�t}��z�83��O����~/j�QX�~)���b�@��b��K2.��U�b`�( +ڮ�{h�%���00�6q���}�>���旑	!s`���\ڽ��L����<W] 2ˊ���q�"r�e����#O��塵4=5�8M�����T��/�'KC�r@ԊV��fh߱��g�U}����a�1��a��)�U��f��ٺ�e`�B�.��S���W�zq�?����V�Z:a��O��>��4�ݹ2q<�^H�jCd����Y��O�5���ɘ'����_E�wZ�z�*z,�������%=��y��6�b�bw��<�s�}�8�q����hN�!>A(wu�����D(����t�!F�?[���>rPu7 +)ߖ>]7�[ӞƳ��&�]������q�e%�>�r�����6z-���<�ǟ���c����ެ^&������U��|@H#�|{��Uji)��Q쓁�׮��G�O�y���W��[lR(+4~ �j6�l��NG(�O�~���c��i,&"���W�\�?��N�B.aC�垕3��U@�!��N�u�)���Bݏl���H��M���5�������!Clr����T��>��A��Z��������g�Դ߈��(V�Q�F��]
�ū:�>�����^4��G͋e���x������aU1�w���B��y����n�qJ'��W�	�`�V	�a!ނ�
K;�]�ۙ��W#����\d��G��K��	6���B@.Q�b�\3w>���[�S��F�jH�P��q�`(�#�P� w�*�c%�"��uIO&wb;��c�m�����<��A�w��3�h%��{&<�ķ͇��2ZB!	�Aڛ����l ����a��Y�T���0O_�j���v4�kp�F�RG�B��_�KOA��;���Rr��L����6%�p6�RwS=�P����X.�~�k�ݱ�^�����#���q[�"��snD���$��+r��3 k<�9�0��lC�C�!
����OA��>�L(	k$?���w��ua����e���(6Yn��Q0��1�$��9��5��_��U�`qs���4���Z��hS� F΢��H�Uyl��z��	Y�=J`
�*���❸Q3��w��\�Y��,�%|x��9t��Q|�� "7P�?y350�۽N�]���Qb�]m���W7�|��&6X|>q�S;��3��Rz�����>1F���hʘ�
�1�"l#CM�|���\��/T�1�T$�YL$�lh,e3��8i����V	��(B�=>��Jv [�
!�?ھ���<�zCJ��l����`��M�Ϲ���#<{�� du�_+�Ho�e�Ym�3�	4k�!d�g�G�U��)(��m�"���c���A�)F^7��?@`�o��%��lS�cfKO�^��F^2`a?�W��K������9V�J�Q����9�`_������՞����͎�57ב3��$��)O㧂'7
O�����d�o��Jb���m�L�o7e�mӺ�h��,5�M���]�}�B(uCVߌ�ʄ]�H_4*r^q�}�U+VJ1_[tӧ����сj�C
x2F�Tdu�N	J�5U�ٳ���O�n�>�X�˯�BxgrS%�ܞ�SU�h�C��G�N���0�&1W_tR���G����W�RR@ ���xʸ�^����#�~�J�yܶ{B���3 ��� ��S�}YuE[8+�C�
�%�@��l�Z�F��<8�wj٬88@�H� ��R�o�	�iǉ�`%H5oɪ+F:���j���oe+���&6ɏ&:����=8ѯ�����p���@g�`�-�_��d�W2rm��� M�+�{w_ES���pBzv`FmF%� �q��F���B�#ct}�׈!T�����7">H�l��_y�;Wh<��Bݹ#�5�dI��#,��27�����m1���x��CZ���S|��ؕ��JD��q�^s���4��@@8���te���d���0�ۦ>�n��{��@"�s�huRpx���#Sහ.�a9���}�M���t�9�D$�O��d����'�����7���A�R���c���5  a�p�eE�o̻�)�)��i�	j�or1B�i����٢�#�O5������{]L�u]�K�C\�J�Qa���Q�("��|@j��扂�u��h(^��J��+(i��d�5�y1/>�#� ����-�f���9}�M��Պ��T�/�)�Z���<ķxf��o/D@X��ΪWi�%�ٞʚ�0��d�^�� s|g�	�D*�xG�k$�c���/����!d�v���lyM�A�^�Nɖ�`M�^���/`U�8����δ�Rx�w���kHӦ @�r�Wp75E�.��p�8��H��/+�U�]L�⠎/c����i��b��`��$:�1� ���Itl9���Hl����#}U�i%Mc�6}�^�k҉#���+dW %�ʭ4P�źd��7��n�_�!���3I���T/٩�p�㭆@��`Ø��?rEI����,��^�e�Mُ�Fa�=yM�������@�hEo��T��T�RE`�48��@��._tAd�^䮑�u-A�[++�㰚H]ƛ%XՇm����V�z�aF$��#�X舤��C�\��<F�hBy^R�op�S_�A�=pfYS��
i� �l�s<��ފ2iJ��t*j\�����)W��C"qUA�@>�Bzw���K.�1|�{ۉ&�������=���$$��U����:�O�Y,��l3�
�s�B1��*~���Y� �Z���f�;D ���7@%t`���y	�,��A�wd�]kz���b�
����'��QȫE�^��pei�{�lb��������;a^��0,�KW��D�#Xe��-�v��T_7F�a ��I(��Y��n�%~�u#�7Q�G��FS=	p���%tP���PH�B��u����n�	�_�-U/��1N���l�apY"N���`�{p�U�^�s�u,p�&��V���&�얔�L�6.^����H�H�n���W��FM.��J[�`?0$I5<���.J�����zפ5U9�(��_��Υ	��B�6��\���A�B�V�<T�V:f�dyzuF�G�3Hq�\�
|���2��q�u��3�}�ǭ{���5F�U� k��������q�*�Q�� �9�w�-�X�MԎ��S{N��4_3�U+Ur23nȿ��pl� ��a�hٕ��̲BRC�e���	�:?m0��vj��r}-��R�W+Q�b�l�5>�:�4�Q�k�e��}���)�r@��̧O�4�y� a��A�j O�PO�ICX���L����m�DXъ	��Z$j_`���s�K�}��uK�8)r�U��v����֋m'w㿷�������OI���*;K�����9�Vl�����9�5�)�����i% W�kq��y��z�zL����B���*�{Xǥ�E-�zS>��n!|qW4ޅ	�M�b��*[����� �Sy����A��>'RgGV�H-q��5�|w?E�A�䭦���-Ћh�7� N�D�"�1_�Tx�Lc.�pk��`���u8�5��*܃P{>H%�d��9��
������t���@��!���+�%'����Α@W�-a~�E��I� ��,_90͝��yHL���#�P�Jm�G`��ɠ�!�_��'�1����1tN��΃C-�@]BW�ٲnVQ%�| ":*��9\?�&]1�!�o�O�K9! gZ�yx���[�a��7�\��cҴ���+)*�^��Ɵ�H2�$r��+T��[څ_؛7W��ި��y��U�}��i�X2/.biq֎�ȷ�!L\�\��K����a����� Q Hf�(F�"z"̽�G�>�]'�P�_����XV�/7�c��
�QgB���Ȇ��9�U�%yz'���1�p�K`5;�ӹpv�����9��6�^Qw66�J̵2�����\5�sP�q��ev�A<,g>M��rK����_��s"�%�Z�j�8���J����˂������.�),����YwR>�`�b�����'٨��ض?XS��wm�/�|���Kܶ��(WI
�ݧ��u|�KX��W2%l����6D��T���ꔼ�i����l�qs?���j��U�T��ݡ���F������,�mA`�ReH�T�� �K�3]حc�T0A��'y���еQ9we�:��/����1�Tmr�'�]<`����v��#�e���(���t"���a7�����dP�[�,�-��|��JXZð1�&�˛�b(Eԁj��Z�È��1ȅ�������N���]���3���[��!e'+���I�;��&5�Ͻ�k��Cϕ<��*��.8D�z<���0t�����\�����z�wjGެ�s�oO��^ˁ�Y�a���B,��8���L����V-S���HU,�!\�R$l����	�ld'�T[F%-I�<#�Ɓ�?D��l���o�d�4e��qe���ݓ]I�T����!"�P�{g,UF���GPg�k��GV>��D���e�EC���-V��Py�$��l-V`�	�C���֢W�O�8����u��R�+���:3]���#*�}�-��n
Bv�7�k�.���'�C�oZ���'@�2��
��M�o�=�jo�$r,z M!�FT�LE��d��r5����g y� 'S��x/Gs��J�1��cn���-8#j&�J$H�����d�/�"Ɯ���$l���su����D}�������s���-=�,Y�������C;K؄4/R�(͙�z&,��U�X|�#�l��Gx-�	�m�_9��$~�],F�gĵW��;s����`�T�ܡ��q�e@�(*�/��-rN���Gl��yh;��Z�46&`5�n����E[�ʔ>��%�P�CE1���0֭ ���'fWHGrNe�r���T�.MjA�ږ�p32���Fi}g��|	�*M�F�M/�ݮu(�Y�1=sH�K�$�Y��<pD������%wYw v�o�/r�O��]�蛷�9�>ī��n7=���xW7U��,��)��iW uP����.��}��Lb����|}Si��_21{ vOli2E�R L �t'cV�P�⡼����T�^����B�WX�;^4�[5�?�tp|7��f���s^���_���}�n���A�����eK�Tz�#\�IMy�8��RR���֝&�c�����P}��e�**��X��!j��m�'z��A���P���b���� ��y�I!"u��� �]#�@x��@zdM̮���~�<o;�K�Z��P���@�n]Y	��K�T�d���ar1�/�̓;����7pBJ�tG+ү�J�-�����E�>�pG��@��O��50Է�H��n�������np��&������xu���/�C,��-�@�w�^�������a��4La�"�R�P}f�}��d"��>�H�l�%@���?��$���+L+!Lk���՚�*s������y�SG����D��b0��q�ځ�cl^�gS̀���:\�,�f�ʞ^��.j�W&��`� ܊Uo�,i�뻪�"�X�^��%�+���[sJO1mm@���Nz!O��l'ӝk-\&��}#�J}���;�ԔB�z�P�����/��A-�LQ��3�Q�D��H��,��\Nf��>q
SkƸp�3�E��`=�W�{����Y�v?��5-�%n8{[���D���L����*�|Ѯr����qG�k�"L�����i�'t�1�=	�Ui�U�HO���~-�O���y�;�.�Lm�(1����8���#hv��+�-�I��l#�^�9��TG��<8��u~��(��y��+C��7�}�����Z�[Ux�{Y}e��My�4�4�,s����D(��p`>��e���.r��x����ni��cL�YfC/\��T�רJe�<v�K�Y�e����X�(B��5C{v>����eD,���N�9L�8��"�U
���ߙB�]�ډ[�:פ�f!��臿qP��F��e8���$��úW ;���m��v�v���4ީ�xL��9e^ r���<�zP���'�x@���ĀT�kԞ7Cȴ�!l�`����$�
�X9�ݸ
 ����T�M�1�9	N�G�ϒ6,�ZD��*شg�`m?zM�� g��$R�Aļ�J�D��M��z</.E����	���g�����x߬�/Ym�8�=|iv��A���Ĕ����ද����@0Ԧ�N�2N�3�Ӊ�J����F^��`�&��p?S"*�g}�e��{�=��>/���x=8�s�'�.^23���`tazJ���{�C]�A$�묷�R)˴�+I�ii����0x)�7,*J�M.}��DTI΀_e�YKH�S��R=t�B����$8uP��[\��UwB$�2�������]�+�Al�W
I��+Ơ�D�~Z�n�)��,D(�f�.���Q]��҄���Ɩ0�)i���ʌ��Tա�w��k+���'`R�O�q{T�yx����|���o�vsk��2�=`Ǐ����[K��u�C߫�rH�e��1��.�-P|@k_v��P�XmߨȦ��-= *~U�J �z��Z{&'�gΕ��ڵ_HZcYoR���8RO{Rd����̾�� �����[�<�}���5�gWJT�b�\g�:y�;���j��i�$2?�.Z0����5��ј�"{��U����x�NMɐ��l�-	X���Bd�J��`����M4�cgK�v�'��y�	���`�6[�i��P�ɡHw9�Z�qv����0�ABc�@/h�/�#u6��F�E3��d˵P���-��j�*������򮏨wY�!O�Xǵ�b�m��~s�&yY��C�f�n+��YGxM���'��2�� qNH�q𪢴��WM��e�DE�lM��.�Xk���a��6ze"e��Z�c}���0�\*;[T���7vh�F�5�h�1͟��@ p�X���(��R�l�Ln�͆�"�n{�4�=M�ji��|�yj�4�5i��;ҡ�	Ey6��Fm���F�=Ff{�&�6	�.�Sr��B����"o.�p9�A-�b�LS��W$�mlp����J��Б�] ��Ҙ��}�""���m�c|�1�]�v�����p��X+�z���r<g~t2��W����F#���gU�����`�l�J;"������ˇ)_�#���m�#?G�0�x%�#��܂^�\Փ�6��:�Tl5s�O,>͏�h����\��fr^��u��fdP	~����XNl"�_WCj�sb#� 2
�*}�!�{��v��8ϓ��)�Y�m �s���~�\{�����7�z:��JЫu����%m-6!Z��h�ٻ����o�N�2BT�����>T�LE	�ŧ��S�,uv홋B��>ga��J�#\C �ܔQ Un��xf�Hǃ���Ac���<�09�M�^�s� tr�/���/2I���`��S5��T4d��q�H���>��ډ�&��v-��eD����9H��D��p�{����I�d�(��ϸd�@�M5��D�E��>,.����p���%�
��q��`?�����z!�u3&����J;sT��/�� �rcv��+��k$M�mdt�"X����sڝ���΍	P8�dn,`��!��w�Y�\�����M�9$���M,"Q>`�iq&�} *���>�r������^���x!������g��b��r���ʶ:�����nX�l���ɚ�u@��sp�9��(��j�m��Ph��L���A���5�����2�߻|5�x������V�����=���O��2oT9���x*��
�!�̵a�@���ǣ��-nu�)�my���o�:Ta�k�<:!��\$�(c��"�����-��:���]��B+fA/Ŭ�|��b�-;�EߚS��}�
܋�<,L�$��cSF3p�]�������`t����zC+4&��
��0.��zf'b���9as"��=����?�8� =.ϰC���XN�v�̏u>�E���/Q���iZ2,C�����l�L�G��X��y�����9�2*3͛���J�'�P�}�W,ls'kZs�̨�[��6�&���FO��۵�D� ͋X_r�n���]�����uR����Ȥ������o��A���k$K�x(�(�;R)Hq󇜐��z��I���К �Rx�Tb/H>��У����p��,;dd�uI�p��~vR�2�N�
�|fA�6�)�2���E�"���7�V��3�&R�V/��������I������ש��W0FA��(Q0�	�%VS�#{��Я\��c+�f�h���$��4���|p�x+Y\��Q��ą���)	��M�oXo����:PqVV��e�8�I��3���@����ӭ���.�`�{���Z����HT�_�3K�N�"R���Y��n�Kq=��9���|�U�k�B�(�5���.��VCY���Jt	W�\�(���A?�V�Q!��0���
n���K�;+m~xl˿����[STn�����J���銮��+�
�O"�SkwTb�`����q3�d�V|�C�F��(��\��:�EF��ڌ����~)������֣g%y�wf�)�O��a�� +���W��x��4��8�[̎�z�(��xJr҃-@-J����d����I��!�l8=H�\������ٺ+�G��Dƭ)���O�T�8b@�[�:�G0CzŔ�gC��5*�n�IYi��/�>p�T4���+�7РY���拰��9�(�wP��\��G����mh.A��/EN�3���	]�x�"sX%?2ʋ���V�`�n�;=p���Y�Lv3sWsc|�<ɱ�r̷�_V�o����_
9k�je�<lM2��&`�����i���L����%�V�Q�~�&�vxkoU4�aDǓ�&���*�ϪV,����zD���c堻��d$]��00�h�`�q!ܺzl���a7�=�Jh_��6
r��$����土���J��Oז�`���ᾡh'�Eq�KD�����~�P��JʓrLQ<[�r���у^����թn<�����^�cT&RT��4����-{��J��ڂ��!!e�Т�KW[#fo7���џ�)�Xq�3���I;r�2��.B�j�)�5�>Wz�c���~X�iYb�Sf����ە����H�Wb��m�5�NgC��M�ꗚu�ZV�����1�{<��"m.��	y��;,}�H�L���!`�BH�qH��ܬ�bH��%G���	���u�l{_��I�Ső��8�D�'J�WjS\R` m����7y������B�ݤ̂����
��i��~���B� ����r��e
�zP���ƾ9��˗%�7j�G0H�������4�B�C3Kr�p�q��ܤQ�3���#46A\�j칥������w!���8�l�V��E��'��� ��E@��F>�&�oe��>	�A�d P�hrЄ�*�@<P�D�Q�rKJ��yɧ���۾����ʤY�7G]M��j�!љ�$�"�>�~����3�;���"���d���y�(�.��	��ZI�A<�A�W+��dro�$b,�wFa�m�"�\��E:�cR%y��R����:'@0�{�SU�TוV۞S]c>�:�<�'�Ǉ	�"�^��8-��><<�2��~&�0��}�Ċ�kG�I�~�8��A�Uqп�V�b���>VD�{�����y1�M��1̸�,��ބ)uJ�;q���߂!�٨�0X[�EGc��[��}�ğ@ɒ���������~�)F�8��\A)���@��ٚ�]���~�yo<�S�)l�M.��	ǯ�b�Q��k�ҵ�J�xcR��L{9F�:�L�g�x�J�1�FFX�����g����vM��A�U|�Jcjl7C<�^o;��_<�hI����9�Ͼ�����-0�J'��	�����������5~ČM�,[`����B[��-����(zH������@�f�Rh,��j�jE��gsN�|(���\.�����z^EY�Q'����C4�\h���8x�r�&#3	H�M��[&(a"�t��}F�`z�_��|�j�نUh����=8�nC�����jy��K�G%��tw��_:P}y�9܊��J
�W��K�8�/:�L�*�� �2{nT����@��m�4̝�H|��Q&�u�qa��p�+l�}����i����[l �P��~sK
ڌ<��56�*��T<�M5 rf-{�@�(�	���);)19%�.<��?��m���VA��L��
~�9���u�B&E��f��4���{4�u^��k���@6i."館*����>������U��H�h����;��m]� �"�a��'i0�  C���Ug��2G�T֟Y2����w�w�����`���ap�M9�b�G��lSvME���գ1?�����	����W�N3��'�I�b,j+:!tڧ�U0zo�O�7	m	c|������л�#ePU2"ULDԆ�Ϧ�R��.z��K{�i�X�|��Ԙ�՞I�@��,k�n3�uÍ��p]��am
�:�aO�$��|~�`�>����%����ПO�~�JPue�O��k�+i�����A��>a���s��:���&�=��`�>*E�di��5֍��: �ܐ����NABw��ê��?'��.�T�.d��;�M�_B��b/8�����E�B��Q8��;�n�b��.��I��eg��l-k��s3��Ñ-U�A�3��W��#sQj[�z�$%��]��X��~졯]�pw $l�k����3Ar��$`u[F?x@��r�f����E=���W���+ͧjMu*�wZ&qZ��uR\���\��y���o���
����vt���+�5Qa�XXǳ����n^5[A�U�ĭ�(��Fe�9���yP�#�X�M�\�!��|���L�3o�`.�������`��LN� ���Z��BG�۳~�c�j�O����꧳�`5��R��FF;?�/�4>��:�����8LW�*Q��Zy,>���*_2nbf�7[�1,�ڐ���/�����[H�k�e�����TK,8Y2q�P�l;��`[�ƶo[h�%�WZ�Xs=JW����n�?�5����]6k0ϱQ�H%
�8�Tt�T�!T� �o�]�kɦ$Z���"��v�����դ��tl�i�I�3�V�*�~�����<���T>a�T`�(��&��,�U��N�l<4A!&"���I�H��nB�#�(�.�x�\���ɩ�#��M��K�]hgw��g�&n�L�j�q1�;��26����v�F��#�xǝ0��|��.�}3�w�tv�4��������X�V�v��=f�ͣ$��<H��ɘ�g�gê��N1�r�w����'m��/���<xѯ=�GJ�%��l�=mǏ�r�+B�:��f���cin�<<�wD%�hl����AeM{�'�J������%��؞@�����ZTrq�M��̠�Ƽ	�-#):CS��aX3��ʊ� ��χit++��K�]�[h�akͽu�sMu��T�}�HD`����㴁P3K�����6YBכ�lk)s@��i<A�Hl`��G��nf�˴p���^�K8\<D��һX�_��
��6�Au�R���yJBKwm�d�p�E���^O��2�����f���:�i�q��D�S�ݪ�#��o>W��֝�nVQF2<��g�w�^?ϵ��"[2��sڏ����$�C���
�$!����.���j�%��qp�j}-�=X΃�i3w��i��l~��iܯ�qr�9��3D'Mr�~��^��ƱC��2��G��A����7���+QI���z�8ܮ ��9�肯�~܈H�=� D����@]�����R!�����˯+|n\�7��ٴ�>�Gx�6�2�蚖܅�t�{����/)~��������{�-]9��b"����_�\l։��~�F|u��̺�ƽ{C�;�t2�������E��O4�cYs��)D�|0�P�3k�8��2�-?!:~����	?"z�����E�EIFlLk#N��WIW%R+���ɪ�9���Ћ?���du��k�TzQ,�t�%�����T~��p�4]�����Ӥ��4ؿ:����1�����w�2�b�`��l6#�`�k'�M/�s"�����c~���[��-����3�j�y��ya6�=9&�m^�pg�]9��U� �1��̎Vq5�7'�7���?i� �D�oeU����W�A.wb�Zv�Y��_��<KA汙�p|���������JĹ!�|+�� (#~�C�}*��1�avNf��$&X�h��V@{�UvX)P�S~j���E8��.;$`�%7Gs�=������[@|3b��������:�!�{�G*Fc!q����<����[�jN�j����� 3�ؔ�w B	�f1����ұס&���cZh�O�6n���䘡�k���K x�jj��/z�SO3��d�Z6�X���f��LN_�5����{��M'"FW�)�������3���|Onl�D��5�/�*�;<W�A���0H]�Lfu��p��@���E7�ߵl�lcj���Wowhc�% �߽�>@�Ie`�+���Ֆr���@��i��bq��hG�<`�J��#�&�̈́�LQ����_\0�XvS�T׊͛h�/�c���}��������HCJ6?,�>!�
�:�♥4"�b�[�L$�����q,�!*�w	�<[=B�r��ĵ[��������.��Nr0Ӹad��;ֶ���Ȼ�i����`Kg#�������F���[jz%_�п�l�%�K5���`�r0"�|���@�&���s��t ��ѷ��ܽ�C�'<���
L��*��i0�RR(49_W
�7y��E�-5�d-K���pf��޻��ń��� ʹ��]ײ������@�-8-*�^�ڄ����Ij��+� +R̀��.�w�;��=bGd\���<����2��+G����e-j6���+�b�3�ߺ�d;~�A�t�T=�I%B;�Z}��?^o���ĭ[�
����q~J�j��.��2�P�O�4�-�ŵf�J��h&������N]��b�%/��)J��8O����j�0�tVn!٣og�r��;*�|�N96܎q��WM�K|�m�R���)�e�%�ks���G� �iG�p��$���=\X�7��n��@�b�G*^!N�h�&��=��us��zs�x����<���3�;A�?�EW��E�!�p�w�c����mu��o|���}ߥ@x�yyu^tnX�6�!�ި�3$�1	9�dl�V=�H�t�]tv�I}'�I\���R{ �S�4y�-
T��5g)J2��v|�`��3 "�C
Fb^���:��������<��\:�֢d�lR8K�P|���'��k���Yn�gN�u�E�0[a�J�D>�o�+������\��ϕ�_��M���IE�k��a�I=�]����J�������DJ��FX�����V��n�?��������#a~
�'R����C$�T�������n�����%T�Z�z�hp�� Եc�А���)�fM�"���QOc��7=yci�l�@kR4ÏW������h�a��K^E�*l	Ձ���Y�=���(�3����8��ᠻQ�Ka���ؤ�FU�C���Zy8��<{�x��A��4�K	��BS
_:c�h�m���sA)�c:������vB�p��Ө�$��*�&BE]pލa�n�б�+�!� !�~y��i��-�� ����DVl>Y�9}>��v�$iBo�Ԁs\B
����R���A�lӅa?[��x�Ǧ{� 5����ϋL���cg_&Ծ�Yˤr_���s��J!G&H�����-���I	ifiw�nL�4p�*$݅x�F�� 8Y� ћ'!p�8
b(�ty��.�a�ݭrG4f�:�u�+����TGl�L<2:x�&��Iׂ�Z]¿e����Ѝ��7H8z�c�T��js'l@%Ộ��e9��HX>so)Y:xw���Oy|��N�cK����)�H��R��Z����m!�9R���g�R��?����n�ֶ@���(��$���: p����-����ldy���MT7��d��X�����Z?r��-c�J7^�A��%�MG�Bd�吜��0�d����F-ڙ"rM�����ǝ���n<r�0V?ZP@���/B(Š;�}`K�	ٍE4h�I�2$����^�ֽ��ir#0�Y�N9�豸��K�0�4R�Yz?[���*���,wR[aΟ�{��D�����C6�/���e�吩��I�I����սظ������!^�����+Gȩyu�
�Y�ӎW� �թH��҅x� �_6EF-̐�+����2j��ݑ]jW�� @��.;�at]����]�d��1  X���d��(��:�Zn0j�d&�^�gأ�lQl�OZ6�h�6��jD�o�V��� ��6b��3���[��S�(F��6g$��f1���c�l�Z�x�$~�ʤ�kA��eȏK��L��M�Pх�.DvSώ��vT/�^M���ք`y(������ĝmt8w�`���2pF�0$ߜ�A���G��4Ȅ{��n�b`� O8��m���9�-U��1�aV]�T����Jh�E���5-2�q�,ю��~�� B^�KoG��n�^���ȇ��6�[b��T�^[�����bx�)�a���u!��^:n�nvt8�vݾ�,��.���X�XVMh,z`���D��9Uۗ�s)��Ǿ΅\���)�d�>���]�Йڌ�hD�g^}��a!�d�I��P�F/ �?����3�>4������dI ��TNKS�Zb�H��!pߔ�[�UF�6V�F/#����@��\�h�>̈́P��j0eV/�n�l�H)�����jT
D&��9��W�����5l���7��s#�''��8
�����[�8��Bշ�?$�~7:D7�O��
�$�,�(�R�M^��~"a4�C7��^^?WDm�i�Lyo��Bե�1ހ](W��n��G�>z��غ��Q��=�u�z�_cG�Z��Y�TT��&����3~�3*"*�ӪNo���~�ܓd���3���2D��)J[�P���H$t������-�R�ءMWl�����c��!g��[/ھ�c��f�e�μ�n���5����TS���^�?�/qRnȨ��_��:�;�.k@�1ѰX�z����^�s��g�}Ir.�+��
)��,Vz�ދ.�
y ���<X���a��������4�u�b�w�c(�b��q䤜}��e"#vJ=�?����np5+<E2眅�Oa-w(�-��F�e�E8���F��]���\��сP�5��r2v�z��5]�)� ��ÅX�%d�u��H��2`���sk
<���=��Fn��8���{�iη1X4�P�7߱-Y�;<��1�>��W��s��/�G��0�9�����v pC(l���^}�)d� ���(j��^0h ������Eq��ZI�;�S���`���[x�@k��C=��ͬ�wp�`=|Aw��o*M~�T�-4�������CQs��>W��^�D�M�@������pTN/�3}�0�8#n.�/�#>+퓚��=�mJ��q��O��Ƌ#Gz�D @��^���'�1p?tS[�.Øg�e�/C���[/�7��ۙ��y��<��/lRw��P_'q6j�Aʾ���f�N����(��xcE���u����p6c�YRI65`'�}�J^�a���o���#�;ɽM�U��o�ρ�H�g}��@ӭ�K|���������`\t����E<C��S	nֿ]0�um��=��Oʂ�uI�l�jg�km�y����k�2T��BC.�(�a'�3�f�������ǟ�6�+ ��m�u�
��GP���@!Sɢo�Z�`�e�%7�͗�F�� ��4V�/���k�.��(��c�Aܲ�!�%8-�ğ�I�,�f��r99PQq�K�8�8�-�A��y�q9<�bJ���Ui�Ty+��
�����/�:������X����$D���MD�4Ԓ��L���#����4��� �Cx���f��n������;���X567#��D�	�.��^�{̏N+�"��9"~�8 b2�:򆢨�W�"��m�����K#TqN�)h9|�me��tE� '��ȱ���J�$��=�����	B��C��d��l/�t9V�Y�6���m����e����o4�>�)�D��~N�rXr��CE	����G��U�j>�cM���ߌS���N牵U�hǿ��N�(�^($��'9vմ���+�xp�T�EV���'GB7�(�*:��1j#f��I�~f�\�L���?^��o#��w��݇��5C����^�X��Ybn��Mߒ��-l|a�2&Y����Z���������i�b�Kd_��`�z4uB#���=?�O�)Q(ۏ��y��:|n�P)bبX�N�h���c�����P�b�U�xN����k��H�H訌5��B�4ZY�
���x��.r$�#���yUt��L���N���*W����7�մ���i���x%�5ִ�3�����z�S��M�3e�|�B�"qCr"r�x�0i����cJ�!�t�r,'w�װ�,�{�\�䒾҇�S�C��I.��`-��g��V]%� �8��=#�|�,m�1���+d���-�D�3�	[ӰӯtE���I;�q(e��]�I�w���M��[�޳mNC����-]Gwg-����'�Eq	
�M4�o����F���97&*�H�Q�'�F9f޵����,�%+��\d��4������"��C�s�~A�ʙJ��.�'m�3�quv9I�/�d?��tuw�����gr��a�U�c�5��;
� r�Y*,bg��i}P��c�4��E�2L�Q8��Em��2�����=#�6�Y$Ǹ�DLc F������Q�EB(b���s��
s���Fj�u���$��&�w�\��J��v�<�����d��$��NCA;�����g�g�����o�ؕ��m�5]z�����v}&~XDLd�p�ٍ����>��&�5�dN$�2��{	LJj��e��+�Ƿ"�4�C���܎!�x��n,N	��Q�0�;0��������[7|�'�<��{竀�<����?�qu1i88�i�i�]#����d�v͢r��n��;�4��!i�[=���C���$��/������߲���b5<�b#����s�+a���� V�+7����PV>˪���-� ,����X��x+�]��v5�>�F�!�g�ͳ�����f���$L����X��)�@֐�AҝβnQ��8U�G����_,�~��[�뗌PzyKF�B�^��`aKKR㱹�2¶�@K�r)� R4��I���t.
�FXB�2���]�9�m:���ִW���)fW���b@	��GO,��	\�=��L���n^o�>sS�����P�w�l$�FD�
����x�vK�T_��u]�#��(��h'�"��~�O�^��n��	Q�T����\��(�@)h!T��(0�s�JUc���>�ʥ�o���Cr(��|d�=��Hc=_�rӮ�*�r;������v`:�ʇ��O�|�6��NPDZ�u�p��|�}C�c��h�-�`�v�1�,t�9ڞ+M�ߛ��Vd�ĬM~ϛ�m]\Ҍ�s-6���5f5�A�#��51�_}�Ϸ%.0���mO������ݢ��w��s�np�Ǖ���"+Ȉ��,}Ļe��DZ��,�^/B�zzJt�??Yv���Z�%mp�OM?�2���}`�_�����Y���!�MR��[2���v�x*�\w�蓗[()b)t��!�����F�x�f"N��l����
��$���PZP'���ȝ~
���c�^�@l����AԤ*b0h��Uݝ:�@,�?�Y�	a����;�2����%�z�Mi=B7��jzf����~�ˎ��nՌ;!dy��>\��R�:��9�^�3[��	Q�7�U(Z�M]�z�KvI�6���  �E2 ���/DA��Z��ʔ���Xc��|�Xfx?Q�@�lǚpHM��|hN<��E[r����X���� �Q�3;��>Ĝ�F��l0�F����lM�A�ֶv��p���|�B�J����S�k����&�0�]Y@�0����|~VG��w�1�s����/�����폪Wǟ	���V]/���9���w����=���=��%q@+��C)ޱ�n�k�Q�8�hA{��� L��_K�7������ÿr��7�zA�J��sX�יr�\<��=��ʤ5U�.D��⢄�c
c�X>��B�;�y����nl�7`�EԿ�(�5o�+XK�!葼���"MDY���DV9}y{�b�����^8_-�>���6�Q+���.��'��p	2��bx�$�E�Z��S�
�E15����d���J��cq��$��Fd���I�+,�)�];ߕh�n�����?���ꠋ�1�&�е!�d�8L��ŉ�xg7�r��7�㛐2���.�=/��r�[�~��>H�@�)����n=6�{4�b��l���}̣����R��EΊ���T�3-e�d�G��xn)C�ܶ��%��.Q5Y�?й���w�[��Ɉ�ښv@=]���P��R���ii:h��#���W�1�/1��b�����VQbG�[�*.A�Ht�0��43����1�tV����H�ڒ���I�Si:'<抩�7l5^6����Jy�O>/���R����9�q�����=@�$�EՂ�s�͡��1���,�t�9���1˄p�A���Os#	������L'{�O�I4��Н�J%\6AV?��Z�0����!�^l��m�8z8����d^�a�BoU�Kh���9���99��*�j�����6VO��fq��{RD���Xdk�6s���Ib��� C�0�>:�%��.N|�R��z'tUM������[��.H�pG܉�����Fu@dހG||M�8���Yq���(��#��Str�J$�;����˒�Mb>?��^DkA�>�����$h����-��3���Xs�>��(���p���a㎧Q��itp-u�RO$S|6y㇬
ٺ,f�1r+1���v<|�/��9��7*�P(���G��FS���G\��X�!��s�E>uʁ.ȩ=�ƕT�v5�OT{]ޞ7@�mJ�U�׌y��֓��Y�ɲ������-��W��FR��O�C����l�S��C�飤fK�\#z=�
KI���䈼
I���e}Q7z��b�v�{c�+ؑ��g��_;�;�z�I�f)�O@Gs�W�+Zu���;�m=TY�2OՇ`Ez�Ű��������1ld��[��I��T�	bd���)�(8�Ebc�a>���[���.R-� X+�n�E0�����1�;_j*dbS����uw�P��O�^a^k�V*A�z�Z������'���\���ā����Ͼ���B<L+�f&�%rs��9�$�q|�|�U��G�ғ#�����e�ƣ6��!,K[�_Z�a��8���'��z�:V8��-M�-ߝս���!��n�J!����톪{��`������Jԩ������Wr���=<���,�w��W��<�H�(5k_� ��/�9DV,p�b�1m/�g;��ھt�d�.�^%T���i�ࡪ~�b�`�r��?�3M@�u�ߕ�����~�Z#�{�tU~�n�L����[�^)�L��#�W��Y�&��^D�zL���m�"p�1�_}=��
(�U9Ln�`Oc�Fҭ�b{�6���[����MI0W���_K�m�y�����'�3r�>���9�,?g�5yi.�<�jض�YJ��@��C>����d ����q/����^3�4�?`��=z�=������յ#�� ����iS�M��>�����|�����~��V� �=���MSl�>C�~��-Ԉ�+ E���# ���"���}�z`�	"�\,�����T�������|�1]��N���!8"�$K�~�(3A��I`II�=1�W�J���R:�+M#��Q��Un.�$��5`t��R��95�D�#�����ĤD���ꃤ�%���猣��Q	W�+`���.~�����{��iͰ��5ȁ�7\�T"׫'+_}}:���� ���@�N�m�a�ڲC�����Q�){E�},W}J7=?=�9�`�t�&q˭@��w�*N9ܱ�&���kd����Rl_�>E��Uj� \�n����=a
]���Z�	�HP���w]'�Po�RK�zH(�{�&�����6��O�?������5�	��L$u�JZ�"������XE�eZ$�E�ƭǄ���*r�1�%R-���7vH1>�	Ooz���[���%w����R��:�HJ�<O�"O����{5�Ȟ��[�
�x��f�V0*(R]��5�㽾�?��w|�K�����Z�8���jQXfa�"�|��m�Ё�C�
�z�����I�?�>��J[�O�v��kИ$�k���yK��zAU��*k|mGeVs M^�S��o��{u�_��k���\��xm6�85�y�= ����f� ؏��>#
�}~\�^��r#k�0{��OC�Y�x1w�MQ:RD�\��������%H#�\2k(�y�k�ҍ:�:}����c���N�-�=�7d �49|};�/������OQə�����YP+k�8b��Ԡpw��8`��7)� x,�,��p	����>��ȇ�?�ɺr*�'����Q��מg�]^�Hv�2�s����^,������p�V?
5��GvQ\Z-��\I,mҗM������Yy�]����
�J�z�}H�L�ܙU���l
����#qJa�HE@��k�]��O?�x���������RU����\�w��?Γn�1j�ppګċ�Z��ֲ�c��S�5�����)�q\�W�ٍ��b}�Yě�5$ʇ�KM������B&z�e/*;1�}������l�LBG��]�D��l��c(ٹ�G9K��6rP�4˞��X<&}ux��[�W����y�e7Ij�{�@E�$�I4����8h�&�-:�z�To[��!�f�0�o���GR���wu����C��� U%��G&Y�`B����0 힢�1��P���s�K.�|�2��zo��ެ��/m��Jf�$ �!��v����7�G|�s��+��9��[2���ǥJ��!d�n��Ή�7lh_�.4=��/�Ё�01x:�z�H�����v�1:�z�%�xHg� A��B��1�l�`�d���̙��m)j	�����;`��'�
��&�������yP��/��xFY�bM�4Wr�-'
�
�pVՃ� ��F4nE�A#L��z;����*װ�������F��}�o�'O��-�d��p9����$��r��٦���f�m�lT�����i�ޜ��9�d*�x�K?%��ꇡ�~��� �����ನ�~�S���x���v���܆A��2��~��_�������V_���f/yωt����aT~-�b1�F��9Q���5=�G`ƙI'0�6�L�
$vҢ��������$A'��<�$8.��"���:�qo��-����=K/QZ�"G*5��u�i����p߲��|̄�B���1�u03@��Z3N嫂i�St��hJe��'�@~��঵�37\���#��.�>�1>��1�a` L���_-��[��XUg�����ʋ7�e  �߭��kb��,�G�Z��8����R�3nY?�������ߦ�v��,v6�4^���1�4���e�������8 ]N�[�W��(�1�*�Ȝ��[kT�Vw(F�B�Ƽ�����ԁ07�~���kk��q�q���ͥh�X���b>8A���A�� �oqf��S�M<��O*W������﫨&�a�J�n�
�S�A���B�o����uE\�<L%�`�7��Ő�3	���I�����b�!�zs�^4��F�j���#z��e�c�_���i�xɵA��6��z���H,O�h�����67��A��Ac�����_nkr��;~�;lt:7"�g�!�$�L��J����&l���^����?B�J���}���;�B�$lo�ܠ�U��|Z(O}6�HY���遆B��j<��a,m?��u"w��Mh� -1�)����.i��M��;���Nq�b� �j3����2�)3����ߜ��0ځ��q5A�*�_Av�!)������(�B�)��)���'�v�:$;��P=�l������HЉ��ҳ���_#�2]X�!�n]�����o��k��ȜQ�>d�g��{�1U�N۟�xgJ8��I�
*�=��u���<Q[�B+��Cga�>��w�?R{�R����T�FS�{�Ay~��v�G�<�{N�	�xL@��ٮ����b?��`�ag3҇����e'�>FYc�0JȐ4�'�Ͳ	W]I4�<�v�5�mh5�����?y�\�F��w��^���6J�ݨz����p��Is�É��'o~3���CZL���z�b��\��P��Zﲟ&	�V�XF�#�8`6��]C�S-��a�u�!m�p��׽}�ܘ�FQ�)��n�,�Gh|�;�D��"�t��������{~�����g�/IE53jF-���)و(���f�+ܤ�g�o�	�����c8Y ��hk�X��Nz��W�]��>���[��6(�v��<�J��U�4wh�E��|VN���N�*���pM��WX�7\+Erx�{��o��2v���	4\7���C�N�X�%�u5S�ɋ"���Q��lp�����9�5�t���y�b��y�=I.K���9I�F� ��or��<,nZ_/]���c��-A�YRi/s؆��>�T�q�E{W��?�%�}����u�C�2a�j��#�Ɵ«�!sɯ!�<�|�hN�ƪ+�sNg2����ğ�C6(b7������*g1%�BG$�;נ����
55�ݪ|�i}��
3>��E~ڿ��ت�� -w
�SF��� n�m�A�Ն�����٢Vbݿ�n"J:��1Uwv�%S ⷕ�� p�_t��C�+�,}���cҮ�{|⑊����Hpf�B����	����)'��f3��ތ�@�9m�m��7)J���G~��@a����!<=��Go�d����B8��nhOAmU�����L0��|b`>�$�1���,$Ťa؟�!��$-�����q4+]�}l7-)"M�N	�	L�k��;��� �8-T'�K5e!��U�bp�����)��}�*��������(򌙀�n~��%�G��PzC�mB� ��({mʁ�J�$�v(z�/���J��3@�!i r��tq �|�n��4O��H��}��V<��҂ggف�g��v����ts�:��J��į���e�,r������E�z1�N���O��`���}<c_�@_sc�hY��=�{ �5��ml�?�K�ʭ�ӶW�ڻ��Br�0B�_��u[�AЬ�+��6o`�UT���@��
p)����v�Tqg��������<'�"s�K&�C�nI��������PO�$>~�gE��
�S�C1��#J3�uM��)�|�3r��q��iT��1��"���X�0��_���Eͳ6|�M�:�I�c�缕��}0�����@���@W%����Id������>i���d$E@��갥��-C�Cf���KU�9���a�?��*yJ�&je�	��& }6_�8bg0���(�[���5-F������M��[�9�G����Y����za���/a�"U&Ô	Tz*D6᲏�#�}l&`'�	�F����6�u3ܪ�v)���2ஏ%<�����ž��ϡ�g����T�`)[s�_�P:j�wWI5�(��T�g�u���y�Y5�V���	w��E�8��'�����H{�֪%,�̓Au
@�pu$B��Փ�;���(�~	�0h�G�Ѣ�D%��ڄ� �ֻ�ݣ�4T�76{�w�4���[]�K��0=9Gڄ�����k1��ʜ��~��X/���� �x�u����v:��ܷ��0Zg�JxF����+�T�N@A�]�%T���XڊeV/�� RԑdzG7�i������}��R�$�a�*����@(.{b�R�����l�Sc!�:�����S��7�P�ce4�]���6ѱ&�/>L�il��+0n32�U���n�����-��dΘ�)��GB8�%`z6sp��ɽwa�� -�yѽѮ�hY�7;88e���,&�� ���)6�~�6^��Ca0R�k�\�:��?��4�����o.@���ۧ���U.Qh*��n��g:ݙ'rm���%dw+�>.9��f��)��AϤ ��{Ɵ���>��WqD3*��f,�=[�G�z�)���bj��H�z��U��=,�b����o�m�Mx̸��g@N�f�C1������WM;-�<M�C�=#�)WN���56��$;�{뤪r��7�&}N��G������6M�p��� ;�# }��+���kD�@��A] �����Y�F�i�`�אJ�h��fT������g`/�`���]���Z��!���V3�2d@�\(��P�o	���#�J����	
�L�SQ��^v���;������0��	���a�O�kkF=k�KG��ؙsL���Q�M Y!ڛLO��J��B�����YE̠>��=�%�d0f޷'G}�+�����;�S�,�ԝ�j��/vA���\��"υeX�2R�6��Uƍ�����A=��B-=��M�1��VR�C�㧋�G�-��g��P����_�!Ghq�#4/И8��@��5sد��!�`)p�}���pj��¾&��A��l��x����B6�(1<����I}��G�Whi$t[���Y�=�B�f&������O��JY���E��v����H��?q��&�Z��7.�Q�PZ��{�*i���|���}�~��X&1^�[G��S��#P�"��?��p��$+[�[=h��+\�L�,D��b>�Ţ�M�L�
��������h��L�9��ٜ���,�%��Bb������=}[�"Ҭ�Č��|�8�x�3�Шr���Ú����������4�Z`��+\��:�|�s�z<����Gt�F�ݏ����lbI٬ˈ1��Y�f�6�sݟ���)рҽL��%</z�6��A�%���gŖ&X�+���˙�᜛���C����>����$E�h�Ҧ-�R;4c�(B�瞞w�Ĺz#ectɞX\����:?^����
�(5Ʌ����qQ��C^�}��$�k�`��B���ٴz4��D����>V��VO�pz�f'��L�(}��1T��Q[��D:��Q(Z�" �5��������"�I�%7�V�z�Q��ż�H���n/��t!��$ρ����yXQ澜���;JXǭɳ�
�����{��Q�sQF�&�k�~\�k>�&��I���N�w�ױ*��fX��r�������!�[�7T��N/��m ���-BM�Ʃ>��~8���_$�}���CwRM���z���iπ���� ?f�X��z#OR�
�y�ٺ��iB�i�Ԕ��H
n�n��`Թ1�6�,7p+�N�?/����L���u�l�'ɥz5�cs�?L�h:�i|6�2��Lt	x��Yx�A{c̱���Y��Y"��L[4wC�نT�B|D�����6��)�+f��v��X�1�5�K����*��-�'Q{Z�v�+�_3��W�b�hϥ!e/�c�]ށ��,Rp� :e�Hyz�6==��q�̺R���P���$[D���s�J7���j��0�?�aq�q�kP�Iے6<3 ����	��O>��\��;��X�Y\���I�A�#x@����^-9��B��X�NfU*�J�{_��,Cj��5��|zE�CRV7N���h�&خ.��KF�ܧ�9���ܞ34}�N�$%�Q�3"��7;��n�K�U��t��3EȈ� eA�_Ee�,��n��u՚E��7����i�PsJ�7�V2���ӄm孋�>J�0/9���2=h���&n�1�sg�����������3gIQ�L0(|gw:�|f����@����M�����_����_E����.wEb{;����"��j��{�?v������a��b�:�S��b����W�*��I�.�>��.:<��{7���<�@G݌M�6�'w@��0$� ��%������i�S���g\4P����""nm´�ȏ68#
��������.2GGs��N�n�o�r�w���%��1�ʄ�W��e����(ɐ'�ݶ�w����~�5,�����'�]Q�r�'�*I�z�C/�ʱH�$��n��_��GaC����(6x���I�ܱI�u֪��2�H�R�~��,Ϯ�e�=Ds�c�p��C�'iv��9�Ly\@������̮x�SpC���"�BM(|�0�ߚFQ!1��3C�<���<J��X��Ę�Ȳ_ũ@
���S|���'��B������,⹴	^�����P���<b�U���_M�w|dC�02�Ϋ���@����oԼ���)Лw��IH�E��m�1.d5;�n��H�������*��|M*B�4م�cӑ؈��� �Y��C%��j��`9���
�C���� �ڃT�Q��e�E��n��p�2�� +�8�����/ =}���N#�_��+Ӡ��� ���"N����4����1�2���_�v<;�a6<�u�� N�Dۣ�,��$|@W�bI�i?:́�U�m)������]��(xyA7P"\��U_��4k��}C���G�e���4�����u��(~y��h�R�BOޙ�qK9F��y�}�s@f�0`�wh����M��\hop����#��ھ��8����dtWޭ�/pM��Q�5�(�c!f�>�,'zP�A��	{��)iU�����x2�մ�U�g_>NI�� ���lX��M.��J���fopm�q=�Ĭ�i��	��h��e�z�v�16&G�&}�>�N���3sV�crf�m}���H �di�6d�^�����ז>����k`Z��q,�:%��\.�vo`��"Aʅw��K��С" �;����'�Pc�R�Kh�m7KmF��[���8�~�VYX��8�l3o��#A¤I�ߨ����7g�>��Ѯ9.Yʱ;��������� �nc�R�(}�)��,���m��5�,@k[y��ǹP8A�t�����C���8-�ufb��1�Z��(��G9��|ȹy���\��_Y�C���ڇT|i%��	G��cH8+�%���rk7��Ŏ��L����y�ź�:M��9}��>�Q���m�&3�]�� *�bm�ב����Q���Ȱ���j���n��v.�(���q��+N�Q/C"�!V'в�#��T��E���Ec�n?��}�D��I��}\.��oq����z���$���C� bv�Ld�q25Ë��R�c=��-���BS�n��H��`^1�HIuP��-H���F��g�[��I�4<��Z/��� 6d�O�>� ���H+
_YSS=z��a��Rw� ���31T�8�&;����sg�+H���Hm<j���0�q+^I
��j��'$�*��Q���權�?FJ1o�`>�'��n;���C�
s���G0�*(����ס`u_�JZg�4IK%���<7�E$ʪi)N���Q{i�޸�;Xq�:<�2x�������vT�o.	��η�� V�F�~0@Y�H��TJmc�����/5����;�)�+آ¤x=ҋ���*\e�U"��j�"��Բ��.�(�s�W�H���I-g$�v���&��&��PsTు
�dUwqO��(����Q�}��z����7E�'cr�ve�@��8���Y]���Y���T>����r����=�/ܐa|ǗPw� �m�+�xrv�/�X>�}S�� ��^��� N��*]����3�G7�f�.��xmѧ�Z�������Ͻ�%^��	�@Pk�Ο <�2�'��!̒�zG���t@`%
��9p
=�
���>�*ڡa�mi6�b �
��{ω��9�?�(�.�%y�?��^��P��qr`
��9�=���l?��ZO�i�@�yΤ�x����,�wIzpz�\��k��y/
��'<$p�W��3��{|��F�T�IwȖh� }�e������L�R�a='p��]qr0>T��yv̩M��l���X䫵pn�\�1�񃗀(F���֖*Ѫ����<c*��H35��������e� 	��:�ڄ���{$� d�l��R�Da���,�7>�q|7lb�K�͈`�*>�츓�,�א	si�0A����eT�"�
���g�OB�4��0�ơ��_v�׬b�0�j�Q$�h��([Gm�� R���O��N~7S��Q-�i21z;�h�,G�d���C�3��;a����g��gƺz�8F�J��G�ݍ� ��� ���"�����1
;r�:P9�~!UX�0�G��$;c�B��ϋH9��~�&,�U��f=�L�?�il�7UmEET<l��
����'����k@����ԭ��jql �D��Ua�V�X|'Ԟ��Xc�D�K'���Rd��GU��8�Y���P��n�J{�qӈ~�~9��<��*�'q�a
 
�kf��M��s�r�w��\M�����P��e�Ғ$[���J���)�]���Q*�+�yY�����&B�z�	T���a��7�ޏ��m��h��{p�&�����a@sO��@P{�L%8۰|���iθ]���˵ �F�V��YԒ�yƽ���P��%[B����ٱ6����?l��li���R�ѫh�k���Xx/v�`5}�S�ޫn�|2>�X�?��Fΐiӯa��x�4��z;'Iga\m݌��i�5ɡ�l��A~�p)����AXy�[Rm�n9���)2	�D6�7:���� )>� ���v�x�w�؜�f�Յ/O��V�������+ov"��f���fvlM�V�'�.��_����8���vz'��yj1óiN?P&�#�$0�PT)�a�����W�`r!�����8>T�ŵ�1����q���|��\T�v�K������|pe?�JĤz��N�T�J$���!����x�J_���H����ZhYΐ�	�@o��^h���:t �^J��T������2��-�io�Es��%�1������{A~L'���sZH������Ϥ?~B����u)�5.%\-H�� �R��<;�Q���	���<
�p�g[8�2��'m�ITR��`���H5�Z8 :��7�71�����?��� �0?È���U�ݹ�SJP�r��V��La��һ����(�*��L�Z�'���9��",C�.�`�x车jq��+�1��{�ٞ�j_ �U�߉�T���7��$��'o���p���>:X�����2(bq�t����cz��?��Ґs$�û�E�b� ��q��K�p�)��*�5\�=l=���#P���_�b�+{���>��O�\���H�T�����ę�9������e��h��T���q?e�v�P�P��L�]��[�pN`D(�}�y�����A�9������x(�P���,�
������EA�O�M$2RQy��x)����'�qY,��l���"��iQ�@�M��$��M�4��3�SP���{1/IB�I$4䇢��l1K/����)����rC���t> �L2��˒�C�|P01�y��U��:�1�f�����QXYG�{e�a�V���e!�<���gc�|���9(�ݨp��ky�cI�V���}Q=��h-��9۲}��E�#���Px�UG&�0�CZfG�ӑ�+�N���� ���IT(��Ƿ�a)b�X��hX�X�	��6��
����qJ���.�-�4ϱ�[ZR�Pٺ
�L� �gp��U,%?UvW�e�;jb��r_M�)�fug&K�uS�����V�g\[�C������,?BJXΩ)�䤂��i#���iY�����#YJn�{���W�W��-,��,��~$q��-�{��˭��P(!���R	����_���}[mR�Fi��}i�g=�'w�M�٩(�$ST�=������?=���F��jȕ{}���ܥ�Ru����J�C��*��Ws�t�%X��Y�0�5b����	��E6�K��)*�&��!�1�#{�5p�/��E�0���Pk�q9��B~V����ȚyV7����Rx���MA%]�a�ʎr��i��y`�* Y6��w@��_f��\n��!V� �)��6+�풃u��;��*T���ͻ���C^����r �t����`�* `a��#���`��Q���k:W�X(?ck��D@}����	t���IJ�^�jE������`-��Xߍ��"k�ᔥ��H||�m�e��|��鞯)%������ �����qQC|�; ݒ���2���8׿��&r�q����ܬ kTY}z4��i�40�9c�`ОȔ��&��ONgy�C�6N5ǇUj()__���m~�Q��|@� e�[���[۳IWisAwg~�
��[� L%H|p|4���2�/r������mL�4���RÕ�l���kzf	��m���дHu\�_�V��t�H	�w�Y�fk E���I�ǣz��(����䖝b���\>�#�����DA51z���E�r�גd�COf��tΦ�8B��S�n<������$�~�y�L�����7�l��\�,�ѫA�a�3")Sl���$>G �lC��R��_:=EdJWZ���2��0�9�����I��3��D�ԟ,/��|������6�t���/`�1������k����������.B-�tf�$\��mX���T�]�~ʕ�l'jS�����+����Y��I���Z�����1�
�B�fZ����+�9y$._����<�BSG�!ԡW�4+R��?����lU��;��N�)�����O�寛�A���?&����|6���6f�-ab�N���U��$��F:�;�����Z�P�<�$~�yWer��b$��=�ĝ�*�J5���uu��`x��_�����7G�Og�Jג槐�����q E˝�� j%�q��J����jzУ��.Bw%6�*�J�;Za��qi?�㈼6�D&ݶ7�β2q�\d�F� �w�6�b �������8�Nj�A:*��cO�O����y ���<.A��Tb�S�(�q:�#e�YQ�<p�!��Sh(}�F�f��hCN`{d��h�2֚�m<�W(�Z�_��ZdC�[O4�n(�U5����tj
<F�v��G�'}+��h�6զ纇�NS�mL��ߦ�@��"�W��g�"uB��SD�m�E*��q�$\�I=�1����[D`\�	��M���W�,��TY��F�i��G���'Y:�a���=���� �~�J�������R��'��+���	J��>��bvJ4��;.Ք�_Wf�|ga��a�;�0���">�x����������|���Y��Ni��ȩj0R��8r�i��,Bg�Vi�l+N<�uh���(�5IX�}lQ��[2;^WE0;!�-�2ߓm��
���c%�Z�=,���fȣ0�,M :��A�w�6Z��8�m�']W��$���ҧ�V��XSZ�MD��î�c�ER#�����*�� � �A����
����9��;��`.���n����d��2��щ��@�ۀc
vWd��>P�S��M	oje�%��91	���o�����Yw�L�^�(�!FTłG����	6���ׁ�$��]��۬�ĜE���L�x�� �( �N�	p�4`_<F��
���G�B�"�\���w�a�~Z|�f��Y"k���ޛJ�}�c9��hR{�5V,�A|�ӧYd�*�}��p`��&�MA#a"P>�kF�8�=�zE��H��D_G9T7o��,�z~a�AE�==<?���k���OĿ����ڨHX�{�mFIҜe[�V�^���m�$Q��{��F܄6�/���a��̆����^�yS�2��V|q��������/�4)�O�,r6Y��t������7�@��D_�4% ����8���9_��p�:��h��j.�ƚfE�@W��h�ǌ9����w@\4Z8����:%��L�s|)��Zd39��i3��-�y�]���A�&{��}�{���{e�AW�_���/2�O���#0_�G�ؗ'�m���ʽ��Rkʃ洋i��uUn;Q���k�Ϊ�'3�EI��g��+S��I8�����̘8�`z	 �@11����+����n�;o�dev�]��f��3G�>��}n��A�$U��=��Xiwe_3]��4�L@�C� ��6�Mٝ��}ؠ�<V��(T�>�-��DI�XG$rtz?o股rN�L3}�����3��׮��u�#NNe�\�t� ��zܓ�A�k�L��፧^G�z����Fo��+F���AF��g%���%i��?1�_��W������ CX8Q�a�������(���("4ObN.��ql^�~� �w���P���
�+`�Wܪ�x/*�no�6ITӗO�tܠ�[8nݝ�$*��D�e���"WfQȲ��%k����$�S�Q��a�*����"�l�]դ���{+�=�n�u���#��"��Tu��6�q-n�F\)\�?��x�^Z�uS��_/< �6�@�p9&pr|�~ܒ��$g&�<���ޒ�-c�K�qS�����������#���b�����	y$D��k-t�2�đ���^Tĩ�����v�2�����������6�i7�W���!8ȝ�#��`�� ��*����~Az�1��Kg薊����ȉ�H~ER�S+Z��� �H����� #r��$VA��q8��X�!�^�S¡�ͮ���3�ґ5�/��!�}��������l��!/ �|®���*�T���-�% "�L�f@���
�|МM�mj2X�Q���`DM����o��cP}���@�0nj�c	�?�}�a��0 \����Mwر9?�K��5��>�(�;��܍��F���<k�j���!�(�6�$:&��c�e<�}�!0e��P�K��@(g�f��*����Hx�.*�%�M~�æ��DWR����c�ww��yp2�{b�%��j	�7�>l%����5̘f�PC��0K�~x�68���M����������V���KCؼR�2֛��e,m�tfp���[��]uV9O7Q�wwB�,p?���~Hڀ�b3E?��d��1��#�e�b����`�? �|�� ߬��q"O.������9��u����xaD�N7#�yU�6�X�<����I�-�
Ȳx�.�H}ҌTt�ub(��]L��.�LV�MU�Z��iŷ����-�7o*��2�@������ C%� ŧ�D|w`3��_���}�޳���t7xU�(����ÖWec}Q3�f��CyY��8�����(1�����a�$C(8}~A����~��@�g`<�����]ʈX"/ I�0|2�� ׁ�m�.ԣW<b4�_��uu�Vb�݋߲��~��i�/j|3"�1���[��ތ�y:T����b�ڨi��g}+h�]D���{�,Z�c��s����hM� �¢�ejEh���r�#| NZ]��u��u��k��a���\S�G�y(���'8h��H.y�����w�G��4�؎��|�8j�P���~���L�=�Cs�>uh����Rs[�{{�C����Ģa��Ĕv��T&�K%������h/�,+����w��.�_J�z��p�5�ĭ�t�^�MGBN���K���E�?g"���<Cu{l�ɶ�q���Tps�GP�`�f���'���2H���Dv���I�C 'r(�Q�|2��"X	�Ӌ�9� �a�`�����MX�Ih~��?�R�Pj�M64���;�DH�d�9�]���ݦr���oiP���R��`A���d̺f�ײ�B��s���|��l)d����b�Q4��'ΉY�<Z�]�϶j�5�˫`�Bz�@zC�)8��p25�-<��2ې],x�b!�����0D��=�����f��G�����y`'��TߤP�X��$Ǩd��I�O�;�����
C(��w[m�N��ci����N��o?ࣴBp�u0Cf�2���Q����Y�X��
���@���D��v�j�dB!\Y	����+�p�,�M$����\5w�����-�y�QK6��N(ԤdAAO��ʻa5J�`�S�KI\���cF�x������� �3J�z�1����8!��Wֈm!�);aU�D��#��9�|>�j��Uu�#���W&3���0y|��6y���eό1�9�6��C8ƚ��o�Ժ~X��Yz�e�^��?��D��tЏ����+T��$���+vY%Q�bQ��X_r�X���R�VM�ݿݨ�AΫ<�a�܆"Ŧ<�B萟�U�c)�UR�g�X�!�<\�e���H����^g�W�R`;@I��2�w#�)<�	��/�[ ���W��#���V��F�w(�M&Cܝ��¢�y�'W��۹� �8�h�a�q
�X��G��	D�;ӟs��������>�����4��+aL�zm�&}S[J��^���u��Vc��8�zd��o=�:�����{�C������7�δ`����"O��dA��0���Y�Ϻ)�fM�L`\�\s]�o�z�p� �g��;�=v��f��M��;ۻ0���JP�|�~�2��O@���v,İ4��������B�ɞ��BRj� �u̷$u�v�'��Q��	a���q��s�w��Ŏ�[+��x�_ztP0��V2Du���ܨ��k���f}ܽ�X�B���4:@G��x��}7h�0�%n�Qd��IC�%5�	�=�E%j6���`WTluU�����Zi�u*)�4+wIa#n�����5y�X+?���#�>�� �٦໦���y��p�!U��l}J�`F"��Ґ����Rsf���&I�uV'BbR^����oW�]'A��B�������}#4�ȧ"o6ޏ��*F�	��rA�+�����M�/|;Gt�6.�K�����pw���1>wn5M���Už�a�ّ����h�|txt�I�B��A�f%�}:�P��0�p�k�fZ��<��� �ɭqŰ��K���20��r�ڬC�+�j`��C� &\���gf,/Tc��}��QƳ�m͈�@�<��ohT��~S#��9�)����W�)����`z�Ј�)�yB����Ri���Q��n9��'�-��ď]v���z*.{�e%b���>?e4� Ņ�[�#���Ċ�i8W�B(����ZjR=��N��G��;Eu�p����4����u�%:�aVjnMJ�.6�IIؼ�2�3�N}�������)πE0NqFԑ,�5�s���~b�������Cp���gV��t���wI3��6ͽ̑j��a��^*D��!|ښ�&e��B7̂Z����u�nD�b��K^��t/��2S��X��O~��J���&qp&̮�����GʉCu���z� 1���y-����]��W�"NN��l���9'�_�����%f���|�q���O~n���/]F�e#�a�̓u|����1chx9JO16Z�\��uI���ӺZ��*�*j�	H��t��rn��Sw�u]}�fA��I��"i��Ģ�9�8}��3o1-D�& p63�_�&*A}�Ȝ ����ڒ��}Iw<$���R����O���/;��r�f�qz����.Ñ^�8r�XJ!�@�f@)Y��3Z��D���耩1:P��o*Y��x��s�I
O�U�}|-v������2�K%��R�k�XUK��㈓�%&b{Ij9[��_l4.�;�.�D܌����|K�/�5��C�<�!~�>3��4�j�x��΍R�{�w���bG�+�C!�^���3���I�R���q2_�f|��-�*�
�Q�s�LvS�օ1B����=��S�e��ITN��Ѱ?w���[pQ��lD�x���F�˖'�|a�S���b�A��Ð����#_�@�w�$l�����։Dg�q�мG2q��R|��_���=���N�K;���l؟<��i,co}֪��i7{�ntCbSpz�������-#����b�^>R��G�P[�З�H\6��������2�~�2y�G�����[69�B����BfH��H#���a�ǣdn0- ��5oą��3S5Rf֒.Y�/��"{0�+�1�Փ�Tn"��j�/ݱTSAb��W��͚�lP�嗉���42��L-�g6͉ە��cn؋-�m�XQ����j��i�5�P-��I��	=����I{��[^��`���r��n��̥B]���7O#��+�����W��>�'�qm���I(���d\L�/�Dl[� �*J��p��t�PA.�j���zbYҡ�'F1ҋ���ͦ-��U�����SUQx�J��R��i��B�<k�9NaW�ً7�T|�M���D��4�8y~�G\��߽��Y~��+n���K�0���6o�v_*L#�`{����t�����B1�\Jވ�V�C(y<ٰ�7�<`f�ޑ��g���U3FfL�����|_r�zuv�Hn���uC�f��'�pƉ���HG�A��Bc�v�s��y���yD,>��~�pI����7�S���Ԅ�֛�$�O���WRk�759���pS� >�n�]�j�	T����U�/R�j�"0dh5�D:��*�cwH�`�ؔ�T ӄ���
=���N����� �JpT��e��qM���q�Ô�\ѥu3���}շ���gl���E8U#��W	>ۿ{�����z��A�����6D�BC��ӱ�#�w/�Um�Ԁy�}@^
e����-��&N�}�|��}'ό�L���bԢ�ҏ�H��U�/A8GA������z���7��"�.ݬ0��M,0MUMRT���d�1㨵6Q ;���~�e#+=�������6��T�$�ё0ٵ��>�0Gc��M�$��	�`L��1��~�`����C�2�v#���ق��>B�{5 o��IJ
=�1���|V�X����H�8���9�a��R��d�2z�K]��/����������J"&q���\���o�8�'�B$��9~B�{F�ǕG���׿�g"]Z �I�2!�I�,`��p�a  ��>�A�4�кf�;D6���AR���J��/0 �?�s�/9���f�|f�c\9���Bk�$�砌��9W�V�7��~
o��$�S��S<��1�=Et&�߾��B�y4j��睃X+(�^|ryv杀ޯO�w �{\Zc��.�In�� �{���X>39}��+�bt���A��&���:Λ�!��<@x��ByvK1�[+��S�޼�R1S�]%�-{��� ��"���/����U��WCg�Q�(�ǥ'?m/�->\1��׺X��;$�$/{�'x�	��DC�� �ʣJP���5#���D;�y�C���2MK=�ʧ<j�=<@n�vd�h��U�-�^K�VS�W���#��_$���l�*~^%�TN1��?'�<$s���%�~I×3���U��p�Q��Y�3h�n ��g1�6H-�!�Q�T_�|ڲ9�Z�G恗�G�u�l�k=�T�)`�hŲ�E�T�x��ȸ��B�����2��.���,Ï��@�� |�_�\�w�2�ep#qQ�vv&��\D���A!2����R`��R�v�f�ksJV
��6:����A5f�s��[�UM�>���uX�4M�ٖٱ�c;�vη6�yg�?l�J�]1���JάN�ls-w|Q�5 ��­��_ iX��eRC�Jj>�(��oJ�����m(�ʞ�������g��@�)���Y[�mq60��T�=H8���0�W���K},������szԯ�X��m�@�`Q�>���q����1
fB��a��/+d&?�g����W8��=��8���\��Ǚ���D�S��Q��b��(���Pw�2"�����?*��^7�9b����n��èh���ά�UKe�AN�z�al�gx��f^A:"Rd��0�O�W^�?E��h)����u��,�~�KU@k\Vk��K�]m)}�^�[+gi�nڅ�U��h v'��J�� m$�n�O�IMR`��ǫ�*u]R�e=�&!A����o��������t���ʞ����ݱ���oy� ��`��%�W�c��G���ۃ8o:�-O��_�N���qqAp��>L8���3,x�l���h1T9CʝĻ{�02��<z2Y��#�K>�K��kOɣα�\��定tKr�x
I�A�fQ�u;�J��x�Ш�^_�I����f����n�@?�vmS07p&=�-nS4�E�=�N�S9���gD�'��F}2��F��EY5�����6���u�G�'��HP��F��8�΄"K�;�)8�]�b�ZN	K���G���S �ݹ����XBʂ��}��g�h?���YXv�Ջ�U'�_�T����͖;c-)9�����؋'#奦��� y�L)=|k������x���0�y{�(,����K���gb��fdBAxD��f�v��C�!���$�ZU�3j�Ic-6#(S���8�*�J"=Tgn=b���}4-�X�vb[N�j��3���A|�J,�U�D+�}�g$��/ @*��;A��"%8����9��)K��/f'؃Fw�3Sh��z w(2�BN�X�/��m5��nX���EĨ��tJ7��+�`��h���V��Rv��&i�� .�z�N���O2�/e���C_ �j:Us�>�K���h��\��s(^R�q2��LYb6lȬbm��)�ȥ,��B�$V�?�c�W{׍��}��Hp�шNa�]��%���Sg&�f�K��|?�bp�M�$W�"�`)���y��8�=���s�/���B�O��!"�EqI����6ɯ��ڀfe�= �$�M�~_AX�I��{��\A:'��8�J��GW�	����?��sy�� ciݩ���Et �3�W'����Wt[:蹝'3��q�]rw���<Pq�2�����ׅN!ך)o�	.`��XE!��1������'�h�x:E�H�wQX���N�>��4/�'阴Pl#�O�!�`W-8X�ܲ��T�U]~y�#H�Vκ��ܯ�b+7j�q��u��z�3�ʽ'���b��J��x[z�HGh &�;�����	�%/D�j��[��\\RkrN��O��e��6Y��;a�J�6Y�#mP��ժ �<�"i�F�"t�t�u7LӰ�cn�&�j�f}U>��Y��9W�i:��D[�/���ǜ�w�D��fv�;�m����`���.�F�KY
�MJJ�<�/~�����6���jL�>5���_�E�P�9�~p5{,!�?�ؕ�� ����%�s	c`J$�Z��� 9����>����r�E����}w��:�un��
����%v^�d���ms{��G��Պy|�a��C�IM�����R �2c�drP+��i�W�z(�?�nN�͑bA5;y�g3�k{z�c~� ��8D�h��8b�~��k����2R:nD�&E9O0fe,��P�>yC|�?},l����ݽ�8�n���};���$v�S�<��'�A���=W�)<�g�F��Ń�>b��Dj�3�FF���J��O�,�l������r�S��f&�5
}�k���&q3�j�]�@�r/AJ&�L��ë��m�tv㌭�Kt������u����$���M��>����lܢ&����E��]��/��W_ �uu z�RgG�3G��3��TC����6�������\�~��$#�ž]X��==LDza,��zǘ��\�?9��v+�#l���_ih���p=��IN �R'6ؑ>	X�N�v[ (Q��ӈ8���Z�@��	8;��<{1��	��Y#��F�9��K�:$@�A�a�d�4T~
(f�C�Տ{Q�Wv��H �Nk�(B�D�T G ����ûm�^����S�嵅�T�)M��W�現�-'KZ��6� �\Qؗ�ɫ���eS˪t>>�w�&�:�M��ek��G�N����;�P�u#vf�@ӌ�T��u�f�Q!Nj���#�s��fP�#�;�󽪮�&��&���Hc��3h��o=��8�|�Pb���e�R ai�#gzm�2����;�˖�"�'�l�;���bq��K+ܝ�Uh�S{����|K��9Q�]��[��L�?YG�6�����RJ��qQu[�*7j�q�4�r<V�����-QN����`�C�l���è"�	!���T�НX���m���KQh`�ܸ8��� ��rq��h�KQ�*
�����GPM_�ff���X�a%��dKOb�^�z����Jh����ngaU�ݩ_ܲ&!5ŝ)���E �as�y�YH��79#_���3@�յ��'����<6�Ǆ��Π֧���|�P� �s�|�;	5)�h��BV~��g���D6�<m�KDj3&a�,��I�ln��HF�����RD6tU �|Y�����g3�@=�����UKY͞���MD!v��vƕ3�e�O2�����s	u�(z�� $��L�<�5Π�AT+�I�AP4F���?��c���U�߭}E��W��(č~�o۽�U��&�߿[B��c��\\7�_�Zk�m6���R,�z�\*��+IT�R�R��Q�>k$cJ$w6����|���{0e�$|�݂�Cy,4d�e?��j����i��G��4;�$xT�Z���w����,�,7�h����GH�>�e�V��#/B�=�!�>>�E�/8�]�-swn3r������1���Té6N$���b�yq� �,f��eIt|�.�_X�V}�:/�V�H*ɺ����+��y�o�'j*	D��Y&���/Ô�E��'���ȋ� =6\��X�uf�K�h���\8�Ã��m%	e�*���؏�<�8"��O�b��cb�[C5�˜|�D(�n����п_ڊ��n`nC5}�Φ$����ͧ��/��a��?4�%�v��K�����	�B0��� � -cM �̸��l��$&~�릨`�5G-� ��))��z����V�!��7Dp���e�v靃jc:�Nw��)�2��:$��	��J����T�u>A�,RX\�O
U6���_Rn�dM�t
r�e��[��{�.M{ �����Zrr��B���|�6̓6dJJ��$�D�[���V5.$��rE�L��%'8�I��5���N�R�Ʃi�����})�e�yIƮ������Yh�_!�fN�Z*�*2�-� �K�0�F�Q�:�R�0r��ȑf�*�}T�@C<�!���9�����fY���)��L�x�KW��o�Q�ߗ*Sm�Q=S��;�fǸ�R�����5�#�����@�!g2��'���80G:Yo�S�'B��lEAea>
�4�Ŋt���ir��˱�F�����S�E[�F� �b�%���y��W�]w���_�^�*P��Gx�đ�WP3�h�������k�@�>�@�gRX׳������q���.C�.�5$�UmB�Ƿ|h��,l�<� �VP3� j��szR�U��R���;)ض���uT�^��S��*_�Jp�	����g¹�b���,������,X.ڔ�~���&!v�t�/E;���Tb���T�]Y,�gex8B3¼0��jx�4ը����v�h�[�^�??��]*ڗ�	�.�^_��%<"�ŀ�%���Zy��`��yLN��a��Cƺ�Dw6�}��`|����5�V=�S�A>���#�Q.�;16����v:�2yudQ�������)Zu��J�^w|&3�%Mv+���sTʧ��h���,�e��:m	V>z�����ppr���Yz�1�+ޜҕ���NQ���
ھ�n������o�����{^�U=��k!��Yh������&�Eś�e��`�%��D�Ѱ�(�g���n7`��!?�O�v�jcp�l���~� �1K�礢1���G�\�U��}��9iКiM]�j��8�o�Ǒ��q��(�T�^�� �2w^s�x"��<���XçD�������\���a�����Z$c�>�I<`�o��%QM��K�P�2��5#?�ܶG櫀Ɋ�ׂ�%^v���ф��v���bw������[���kV �_LG	�'J9���ϣ�Ħc�\�j��P���8�VK��]��C(/���D{�ŗ�$>�<����=G�b'"��ɺ�Hq�w�I�E%ť���e��>5mS��6��Rt�G;���
z��ojP_6	`MY`��i�u?ѧ����
����:��/��v`���iω������\��ݝ����FG�ϧ�!�{�:g�7yE��C �/5�����(k\-aw��i]� ���*q�XT��Y�'�s[E$b{��b�c��1<�S���jG�:4���Bk%��f�1�><�lM� u�{�}�����|�&�G��+�S�u5/�S	�g��� _�{�-"�~��i氝�Z�����������T�Z��͛����nU��3oG!���l'Rs�3�S���fB���q��٬������t�[&�
wd��܌�U�cB�ljJ�N�J�cϋkr%5���{��Zi� V�#MqǵG.����A��7�+V�t)Y��¸�@�,ø��q��3�]�����O+K^��Hj�M��-�<h�����[k�����Q��}�x%-d|��{&�y1b�[�~Œ�i�<�&��Z��ȍv����q����,Z�^�h�!(摂�LȐM�_��\1�bf���s].QI�v�Ҁ���S���W�?	F	�W����]�Eܠ�<�8�W��|���کa�m0����&�����ey����m�M�z-���N)�����Lu����m}�����f5���,0б��⿧�V�9�E9�˚����g��_�_�r���q4�� ���	]���	�0��v�-׭l&u�������_?s`V��A~h>]���gk�_ݪSQ��F��`g� azT�p�=#n��H�p6׏��jnhP�fܺOS4{��0X���>�u����O�ӌ�1��8�M�^�J$��(P�7�M6��$oe��9yx�z[���5ulHp�:������'p ϦeP��P���+��\�O��w�<�Q%�m�v�b R	���34��l6��;z~�<������6ү�w&Հ���Y?�=��2Q���}"�s��T+)��-C��!��&j΍�ݲ1��~�?1`������îS aXYH4�Y�ƕj| ��	�y�Q�Q�i�B�E��o��\��`�]qk�jb�^��&BT��rpT��L?`?���,��� xU�}����
D1��{��m��N�>�,F���%
��#A��6)��U����n��d0��v�$������㏒�g[�� UD�Te}W�Ϋ�D�7G�׊��2����^~�������[<�7�~k�j�S�N$���t�6���]�rbF	��D [�.�a��G񔙑Nþ�ɻv�F���6��p|�*�߲rM��@	kƒ�dIH��� zņ�F��g�0�j���H��#X=�)��o�@^g�'=\#��-1����ό�:[��U-<�Q��h��^�
gr��ŕ��'��(��Ҏ�77�	�|�(��������n,߶��<�&wb�ضkt�c�N����`�Jd��-����e��u�bGc�2P�>t�L�{���UT��[1�c�\�,�C2�Pc%��
�0%�I��Fڛ9���;��ĵ,W2��q
Y�Hf�;��,��x9�h���������UP����\�&,J�m$�w�_dѻu@���e�b���[�*Sڀ���
��_�Ew�3$�6i�R�Mlm��sˮ_�F�M\3Ɏ `�QM�(c�*p��Lm��h|h�TX#fc�ܭ��h�4��|b+h��ܢO�m�xr������E�H{��-��˩�^�|-% &de~TI�Ք,�fh�ƻ0�,3���>�-�����N���-��#
҄JN_��ɦ�-]R��gJ�s��PJmS�g��a�ԗ.���ʯ�/��3��*���}VZ��cr����-�������vb����ڰψJ�H�ǕB
Ÿ,�ɰv"��v`�,���^�7H�Q��I�����4mq����|�f;�kդ5_����|�F���ßJ�1��0�o��6�jGAD����<�G�h-���9cJ6��x�n�GK��--Y��2���3��X��e����7{�/Ĕ��fR��a���察!��â�����1���;�ʪ��r�h�9�x_�>�
~�BqG�}�}P��&��i_��"�bn��b�W��(�Tr��<@$����qD/ď���o	O���̼�5=�ޜ�e����;�h�J��
�J3�PK�'�҄�zg�o�q��N��4��HiA�?sf~Ѩ���?1������(�7-^�u� ���?��֥I��%�ձ�.�jyz�K4�Z��ؐ��uz�;&,��ξ�8�I߯X$.���{n��N�v5Q�H���s���m�*�����㭸2dW����#��/���:)���O��Xk�`���r�.���^x2Ω��7��"��v��4
�ݝ$IЛ=����t��%���V�~����M�Ŋ�ή��$5 �d!P�U/�Q���3�n� �;����ϖێ�а�/hbN �5�Na%�u�^�e��i�E�B����=�A�����D�3�@{f�?1� ���egu��̓̐CeĤ{;�04����-�v��%��n2��:r���iU���iB7A��q> +
�$V�o���� 9N�"��D&��:��j��yBŦR�����0u^��$�<��gә�o�)�]��6���m1U�g�;�锋�X̍��t�.�%ä�N �+X1c��X޷�0"�(�c��84���pT�.��Ӵ�o+��I��iRF���hu���u�A����rH<�M̺8�a����3��?`�ݡi��5�{J{�u�L_�V�u�o�.l����]]�r���Jӭ �zC��C�2:��1'������]tan�J�8���z#_�[{���%����xe�:`?�W?�]_���z�4�z-+�j�8���mxX�I*�Ӈ�P;����,��5k���ֶ |��*]�|S�~�+Vj�pU�2-9��Xj% X�18��gq��x\d���ڌ�Uwy�D�,!.dfiu��C8������
�SEP���@Y��kM�]�N�qU����߉^�.�o����J�U_�SK	C���M|0�}�iH�
C�Or�I�������Gd3�����1��l(�u�g<�?T%<�E	���-Ox�,�.ᤧ`P���ј�����!��B��@��"��|G��	�f4�)~5���'�a~Ԭ�b�+�|�mȆ�@q[���Eӊ�b4I!�"^�!{�f���X#l{����/��-PL�b�FY��j����li�{�7�n��('mtQ�ۣ=��k?�Zoٚ��D8���R��ݖf�JtX�'�r�,\>m䑟�	����ޱ�{X����q�c�[��M��{l<�:�&�nJP���'c�Ic��+���u�C�c�k�Ly,@`=*O�t�Q�&`P=0�7r�V�y�Z=�2^�9��Kiq����g&DP��gq��&�3>g��M�:��B� ���b��6�.��@��[�;�b	��N���8�L�m�h����CAj��� 4�||,�R(�K�c�f��9z�}0���t�����l�+�� ��!��t��v �x�����,����S�Ƹ��v9c�k|+����[���n�2��>$gڌ���E�5�.��G=��Ԋ��ξ�1-����r�`^s0=�WM�������&���4zE	d��UX�'C$i��� �XB�D�@�b��]���0�?3��hX��q�Ǔ�lk�E)��UQ)p�c�s1�6��ql�t����q�c
rfG�Wu�a���1��O�Pu���X���my`~u/��z<TV��$��� �,O|�d�%�2O�u*M��P%�m���1�V���~����c��O(����mC����T���}
���K��b8��1�X�oA�xU��zl��Q��۳����<���9{��Tϐ��ЇLy_�韌��c��C�v�'�I�Y8{U$���x*@a��X�W��H'���_���o��{T5<�� HF��S�U:I<		C?f�/c���ui�����$*i�qjūTۜO�!Q���Z��5�!��~%��"X;���)�*��s�2�%�lEO+ ���^4��,om�Zm�ע͎�?�,�Ev�9A��8"ݺ��a�寢����1v�����ǣȭ#F��S�p⒏Rb�"�&�y��\31x��M������d����u0:8��{|���`-Y���^�6z�T��ۋ��i��Qĭ�u36�-�,�/����;Ӱ��7���μ�@剴|'�j�[��z��R���:ޙ���+X�!
�C�@������!�~�L@Q�_�G7'qO��ͨ|�ϛ�L.��f'�������(�r�k<���M�V���˒DW<t��0�l5�����g��&=-".�"8��ŋ�	�w��j��I���Q% k� (��}Ej�߾��<�
��o��^~;��7n��M-��<N�	P�T*U�y[�|�b6a���%�i�[Un�f�g}��N�r�=:��}�|CS�H%`�j��K�5_�#�2�]U�c�S�� ��V.���_۠�$Ŏ�2ء�m_�j�3�+ht�!5Է�[[�X%��؍v^^��s�hȰ�B������\��I��cĽzk����	�5�����M�d�(��s�H�|����Q���DS�����0��G8y2Ӵ��nz�bb��s+��� ����w�ԷƂ-�<��Q��)�Zg�[��O�Ν��қ�j��}¡�7B��&�Ɖ�u�@a�W���i�Hh&E�@E�k7_֎�t��G"�`�+�6��X:�4U|�gFH��d�q�£�
R�(�X>T�	@��>�>$�I���*�GA����@��H}�M�x4��
H䓬 �L&�ԍ�I�k[��h��fYA��3'���3f 8�6W�;��Ʊ! RjF\L�W�Ϳcia�����tޝc?�囜�Yr��4;�L�%�V�a�	���1�5�f�h8��	�SZI0~��j5փn�`��|�H�=^�e�/1':��	�m1�TǒAڭhm�8����˺�x�����,H�n9ŉ�.>oTD�~�P0�?;%�_q��K�𥒖�7�k�����a{L���
��s�� ���q ��J�v���Cl��v(������d�� �}�TY1P6.d$i�oe�m��.*^jǇ6M����d0����6�6�óԌ��^�N3�H��U�h���3�}@��@?���bϽ��l�/h@G��(?`bX��;HKVd&�4�t0�b�g%ٱ�)9L5��=� ;<���3�]!�.�sdi���L�ȏ��Z9(�@��n�R�l�X-��1IҰ��Д���_k�T
 ꚧ��BڤM�?��vB[��v��)n���{�ݲ7UG�l4�+s?���LbÓ�����Q��"AIBt�=��V�����s[��}E)��O1۟�S$MdX���i�8� ��8��75��ؗ��G!?��+�1	�ލ]��u���};���\���˘�i]N�#����~���}ɛp�<#���µ����T� �W��[�g�Q��+�����k����Ij*�Q{9�"K.oL��������r<�L�|Mf�o޲�]G���lC�\�2:���q�`4�&��(����ς�#�h�lO�m��b�=�3�[�7q�a�d��R��_2_9jp�IFd�#:��6dƴ2�	;�y�G�)�Bo����m!��&,�
� �oNE���1��K�ta��(��� 6��$>s���8��@@��Z8���o{G�(�K�j�5^|?-�-8���a8\���L#)o��k1�䯬�;�����T�{BT@���6�$zu)ؚQk��Oc�[��Mn��t#]SV6��k���%��j�p�/Ϊ�M?�O�egejC���T��Fx��m�4��m��� V[��`U��:�=���x�Ft2�N���K!�8���n�in�K��{���L~@d}\\b%�g�K����U�O�k��\N#b�E�!��o�[DZ��i�`Az^�м͓�P��5��:�;<��$�A�@�`����ܬf���(\����b-�RS��6F���sh��#��J� �vM�V:d6�Ab&qI��AMpl	V��!��^c>4|���2[�����q�1�ykoը���\H�$j�h��v�LZq���1%�E#ܟ��������Of�=���:��Hf�ϵ��Y��nb�g��s���N��u�nB���zM(n�P��p?.JV�X{A�ՠ�`�h\�@d���M4��j���Q";{F1�)q���GT$(O��z7�ڽ�8y�><����Ǻ~)&����m����H�V9��p���&:��(՝����h�W�����m�>N�({K��!�\�����J���kI`�+Ȋ}v��B8�eJ��6��]�p��Đ������+�P�@e8.4^G�y�W���r~�+��y��� �<�y�e��j��O�;�&Sg��a?l]��F�Zdno�{㲵�;�H�p�ە�?�zL0K��J��g�]��*ԛ=U�X=�^4/kF�*N�Gn����q���>sF���`�-~±��4�G��}�m��94>�R�����$�%wӜ!��7�`���ȑ��/qNM�|���D.%B�`�Q�߻��`�]���'3��]�'��%�Z��}b�5�����}�~
���G�-Mţi|ai�!0�ٮ-��!$	t��כW�j ��- �[��`~pRmwY�wI|i�����%�	�^��)����z�ryK�;-��7^��e9P;m�^/�s����'{R�d�{M g���[�I:E�6�hF�@��3`yx��Տ�Q�JŶ�<��G*���Uv@#h�&�@���y�%	�B�6A�{�$y3���[���y�u@I'�LM��tɕ�� �M�G��m�a���pdC}��Q�:.|��B��L�~�X�D�U��0p=xb�c�J�#熕�Ɏ-8OC*�Aܸ'LqXb���S��6)������������R�3'�G,y�(>�z�0ew{lh̀_w8([�J��R$�})���*�ݐH���]γ�e�_��5̸`�����@�sT�-����T|?��н���3/��?�h�kK�%p[���^C/iP'E3�j:"���>�̻
�̈����D-�/��c�U���o�߹��4��6�R��kr��/+)=qq!�ŏ o���>��[��l��,B*�M�N?=oIߚ�W!k����U�.�������>�p�Y8��*B#gO2h[u�yV��ر؏ˋvv�n:��Ћ��.�X�g�2y��%f��4�%�����zP�+���y
k/��[�d{U���?��9���j莴�ؤé�
\��w�r�1_�[m��_'��ʈ$=S(������JN�:��У���������Ic<po8Myu�^�45"�h���۸�wP�ۧ�>gp3nAa4��jj�0F�Sh��U�S��q*S�Ĝ�	zy�ϯ�t���g~��tl_�����c��F���L>�8�r��^�ޫ�u�z&�)������aVȶ�j-����U|��i�F��O��V,��hbv���*������
q��M8k9ɶ��h���?�ހ�3�Z�/�K�����`۷�S2$�.�jJCM9����Do�YA73O�k�"U�x�Z����G��k���2���&`/üH�x�Cp
w��Od�Cp���|#��Pq��� ^t��v޻t��%*=�O���?�Ēn �G2hY��4�����[Uh��e�J��n�h�
�S��&��]ӯ3<�%�_�`֥���|��R���ue�j���ٔ�I�����
���M{��|�1��'�� �:��U�@�v4��ܼ!/���#�s�a4+��q͝�	3H����U�$L�	j93啡�����]I(���� ��17��?%I"�L�[M��a��h�u��Q��9��n	L�Rz��y�,��ß��YB�+('��|*j���
��7�E������{�KZ&h�?��8)f�G��ߏ�ϊ|��+������o!�˴T�d��ϫ=���h���i�e��oW�=$Y��]�p0�ru�6Hiq�2�o�L��Sn�UyEw��	=���;��G��3�l��<�����$@�kk�����c���F�H\D����g�p����9ՌJVJܕp����(��yP8��^_���U�{��hK�x[@T�Ш2,W6hee�U,#PG�f�6>��V�]�M3ת>�O"����Ƕ�������U-?�/��=j������e%|������ő�m�tNkB[���]t��7��5Ǡ�5=n����O���<R{P��VnǮw�l�rJ�I-圆қ��:�M���V���iB��Ä���A��p�
��_�o���S��V��'�̋ ��BV�*0������8�V�*@��N�릝��W��RC�� ���/�l�2�����R��Ob-A���)긄pK�\����r���q:SM�N�E�)cu�+!}�R�4�̕g>�^�Գ��Sl�o�T�upKk���u*�r?��L��,+��e�{kJ���)��]��rid��A5��]�|�����?���g�@  �?f��9����(����QH�NOC1���$���J-��Q���AcܔQ�nw5So���	��Z�!�[��A { Ӱ^w��ǚ�OB\�C��-ċ�� s��%hW�D� ��4�j��uɎt�����x"eJ�����7�r��u���H�z+k(>R�k��]�>Q�Ÿ�i���Y��#3k:�Ҕ7��#��<c��h���]WN��o�p�C��z��"d��,�Y�E��H-�/��l�R�M�[�@m���x�a�_�H�/J�auy5o�(7���O)�CsJa�x��������:X8�<LD�?��ʥ�Z��R��h@�u��4B�\��`�#�hU���W<�^d����q�x� ~�-�[��8L,��^�ܵ�~&D��Nt:�XnȪ �]}f����0���>�FR�Q6���E���i��L0����� ���$��7"�>����$f�����͛��/6�{�g����Ф�i��:��Հ�՗)���1
/�!5��Dd�H��ZE2�dVg���"hyJ%0���N�o8/�Z�]e;�?0z^]�n�[���5����W��ΌHs}�!���Dcv0ơ�O�e�܂��*�(�u��K:m�J�4���K�����TIf��fG0`P�L���t�<Yb�x����vU�q�� ����c�-t?�C��Iw1:�g}�u.'��yS����9��+'�@{0V��}";�ٽ}�_(��qת�����f_�\��R�4c`��i8����g���D�@9
��u�2"����8=��'qڛ@
ƾV�>��[�� ���m��z��P�� ��z��aj���~t傗qwE?�|l��Z��N�čK}��덭�ݐ�(38�&?�HyP@Yi��ۀLGq}��4c�q��W7Y��F���<���s3*�p��AC�.d�F� �@��sn�
G���;zj\[1ѫ�Cv\�<�)�u���AM��y^6�%��7�8R�ǳ R����GƤ�/w����݊��9�k������[a1c���
 �2��q��f�0����F�k����}~��{�Ii���ʌi��i�;�t��t	E�Dr���z�E`���=c�p�3�c��7�{��`��,~�]Mc�$��ҁ�\Q����Z&g�꼱s�A��U0f���P1�I��;�^(� v��В����;	�ha���!���@=Ys��њ|�R/��g:w9dQ'�pa�Lv��!�	ʕ\��@?j�F�R���}i����cB�Ga���w�-�s��A�GΊ�L"QK1������
+JrМk��hR���>O�3�e�`�S
|]��п@��F'1�Xh:@a�#�%wB�D�nQqg��u�r\߷>��T,z�  ��h_]Ϯ���K�������S+X��Ab7t�`�t�S��R�Jj~5�����giN�\̠UE��� �
��s�M#
��0��+5��
�@~)Jk��o�S�-�i('	�kH����^�42��JAut@��`Ҏ*�+�mb+*bJ�ĈN�K�"f�Ũ=S��',��h��@�c�H~S�*�0��{�Z��4�|�n�9-n00<%�:�8����'̫;A~8v�%��r�C��O2ap��K ��}�����`����x�¢���y�.5Aag�l��.Ӹ }u;�K�oun�\�)�Z��e2k:RS�H~���~��G!����+[8���?Af"��'POzp�O��N�B�n$��(֡��"��;�gHW5FA胚�^�r$�f�|�Mu����S��'�y�
e�:���(��l m�������b�x�!�!x����{���,��6��`���w0�Q�Mw�\<��B'Ė{j����S4	F�5�p�P�u��&�zӭ�����Y��ڄq�ōC`����nA�JspX���%�tS�$K�,�Ė8L��c��Ҷ��*;�aD]�n�!����5�7� q�#k#!��G5��V�4��C��]���~�7ĥd�Bn�k	��t��b��ƹ�Y<15|k)w�UƘnҫ���[6qQ��T��Z-����q�&�5��N��a�I�T��)����||~P�?B��p�_�BO9���#�b�9hG䐮)7�\����222���[�+�T&���W�¯��9��fN�(5!aݬ��(��|�SV@z��\���	��pD��I�N�Q�C��R!�>�����G<|Ľ����?��=72��w�>X�=VD�V�qcύ)���;!�Q��w8M��ݙ�2�ﴹ���}y��#�:�X�-�W�F!�9���B60Mv�PjX�q��&�GDg���M�k���\V���������4fu� �i�s�.&��t�/Zu`\a�$��u�����2y?H��L��B�v\�.l�55�Cpx�$��=y
�	Ӳ�i�^+]����V��'��͵O�~������H��k_'��6_�x7��$ԭ�u@���a��.6�VkJ����{3Y��{���{��-s��;�	��/��h�	��!�X�80���el���\�QZ�d�Kq�'S��^�$�|̥����Y������s*�ټUKJ����*��H�f����[�m<J<���=&�Q�R��tLF���èk1��m*�d��x����%�V���P�K<!�Sv��)/�7�&��P%�^�YeĪN���|4q)x~�_j��|�f`c��Ղ"~�=0��{�8�/�
 t>bܖлY��<\�����iA����6Z����3'A� X#�t��A'�!�0<
o�{S�0�:/U�(�F�ⱱl��Н­@�G^m>�|��)K{A��g1c�!�{/4'fv�~��1��ܰ|vH�#wͳ�����������ك��'��b{��m��۬�� �W�!�=M%��xR�n=[�@Σ��J�<ѡ��Pқ�gN�QH�s�6��_[�/�~�)Or�>as��wq��jW�[�J�L$9�܇Q�^yH��b��D�(lR:R^�bCD#�oٳ��w�h
o����C75R��TM���5� /*arh�?;`i���w�)}>�"`��+��A�82����Xb��DCq�gpŲ��i��"�m}�(e
�e�BJ*�=����!��pp��`%��]:��Ԟw� ���x"����Hi,�J/����kb)�
��lv�m��0F�;> `H9k�VJM�M��8r��@F势��J
�;�Y�^�@���L��B���ƟKkjn\:�lӄk��v=�\�μ������q��A+�~���V�{R����k�^��-��e���L���I=$����V�3r}���U�x��¦I�\`����3�K�8Q�=�0Kz�ڔ���J�����������2�ڟ�/},�z��g�+G��Pe�6�P���ː{4�D��Q�L�,zQ,���{yu����d8b����\"��n}%�U��!��K����V4��x�8$\�J�bQB\�|[���KuBË\�L'U͖��M' �\[ھ��5<U��������e:�P�Tm���=�D��j�փ�G#�����8���k��<�b}[}�����[�^�]�`�^6RJ�Ê�On���`P^��� ����m��6�����0K��uQ�����rN2`��_@�w����E<5j���ڟ,�Ym��#���P$G��2��e��M�]���G}���	M[����zv��+/��������M<X]��{���G����T���?�ea�K'�YQ���=2sd1��!y�d���^�fx��P���#?��pG���Y�Ɠ�i~��s�]EP<�Y�cO�������q0ò�ďVJ-_�"Qg��dG�j�p�/?�g5$���F��� /EvV�$8�:��o&P�͘)^�&����P���ϋ�މ�^�ΆDn��\�k����q�+ ���/%����vK�M��z[�z+q�%��`�{�7���n�Q�Ic�.��9�2u��.w�MHv_�-z5A��R����=x�Aħ��h�+��Ɲ�+���\ڴU���-�����b��0{e�q��2a�#_�����_#9l����D!��������o��f's���_������}�zߒB����5�!_.�Ag�P\m2� �y;��A�L� & �FU 1Z�Է�m\�O��y#6z
��m�s43JM�-R��>I<q%�}�8!�]��:^	D:��n�<)�KM^�+]����ڬ�Ӷ��2��{'|Z��)搘��לk�7�)�鎃8�[����a��,�M�#$Q[�JAO��kyJ@2}�� X�u9�NI�>;岅v;e�]�J�.��b5G���I�&�G�]��O��j@Ӑum:��u��xy��Ƚ��p��M���?�R����f,�Y5v��4e����v\E8���^��a�!�lΰ)n��>A��׺�T���Q����86�i�i�gC]��L�z���� @���D9�Y�`o2Ǫ���ؠ+�*�t�l��b�jxm(���� ��4�a}�V_�@�|��=���^8�P����Y^����{�`H᷉��E_^豼�y�J�ڰ�q�!('�>��ݿQ��t���< ���c�#�U�1�����bE��XR&/|�%Wڔ��Ҷd腴��c
Љ��z�����O0?TNr��I�FL�a���.A�tS\ª�����
�i��!��.�N)o���G�� ���f���0�ϵ���"�����?�
&d����.�kul�js9?�����cX���&k��\���P-���,�v��Szn_��XQ@�f�.-XB�uA�9I�6��7���X���E���֖p!RT��_��<ZYϙ�9�Kc�,�<�N��M����M:�ϔ��KfT���m�>3!1t�z�i����;�K׳A��gI��a�����]@¤�_e��8`%4e���u֓�$�q�M���������4s������2���m*�v �Wr/���6�Z��d�*q��h��6	)����D�����{�q	 �9׿���������}�? ~@��L�O�E�Հ8�7�h��"��+�C��x&	}�o��U?�M�ٲœMW/����(wZd��}Q��4�e- �y�Kt%����}���wi?�����0��Z�[�p�E��雃��w��>i�@W{r�c��L�=���S�v٪��"�Я��1� -�ȯܿ����e����3z�O'�_��T�\<��.^GC4�Y(�)b�ڭ��{Z0�k��G���/��;eՂ�}�����p����2b|;�����R�(h[z���sļk�\�k��4�Q��K�3ܔc��V��m�kf�#��UXN�3l����6���`���k����;��d�=�s���_~�h
�Ua�dhp�H�,�=,�����q1�z���;�+
R�6�p��S$'�-B�Ghx�V^h��F��a��!�6�9"�ZW-�j1�	L�C����qW��i0�T>,��Ϸ�"].I@�}��C"*n4���|���@#3�����n��9q���K�Ǚc� F��볒���-S��&���#����� �a��2q�Ǆ4�f�V�ZVr�x5Nq�l3��������Dڪ�� J��y�^`�kZ Q�.9
[$h�Z��Jrw,Vw}s#��߭&�Ql@\�o=��E^�$9ک��e�~��Z �c�nl�+C�~#kd�_݅�W��L���T�!�й|�A)sΜ�>>�ԋn�&�WW�M��搉�g��P��o�u�q%�x�p�Ƭ����YQֻPO��t�����z�;xo���QO�LP�e�e��"!Z�w��`Ջjs�_��W�G�6d;Y�3 �: �\]F�M�M�8�� p�����A9D��z�����U$C�.�����; ��C��!^�(��襀8{b��e��9RvGs|F��=��DX�ě��r]'*wG�j�����͂�"r��S%�9�ʉQ/����:P�ye�\ �I�;0:�$�/��wPJH~��H K����$XAAi
�)������3�s�l�R4�!��l�Վ@��������:�t��\�s�C
yf6J�9F�1HޗaN�+Z{�F/)��^/����`? ��[������˨b~9[��L\�Jg����+:XB��3�h�֘8�y9�O3����>�o]3y�v��� �hV.6B鋠�ے�H�sw�0�^�����x����Vu0�&c>�:�q4&T�z�L�E�<@��GD�Zy;�ʺ���P��$�H���4݉ �и,�N�2j��E�=l�
��j���?mT~�R���
��in���'�#���%��2�D��	"{/|
���~��K�T(r��{"�#�$��L��;)Kd�>�xo���j�i�c�^�M1�
�M=� 8|p���&~$5
�b�����4;<�şX���8�R-;)E���B�[�ϵ�o��r'm=gj�ak��
���Zu�r���pU��Eg�-}i �^%�5 x6)���~0��C���}F���o����yM�n���V��D�#�%_"=�h�E�.��L�hsv�-��M�8���T�,�����{� �'!�"�G� =1&3�&����wlms��,�D1�~���J��1P�V���&+��|�Y�g��wr6��$p���#7�,�V���l\��dz����n+z���{��1]6�dV�7�f&����h��+l��*AKˆ���O����)R���%?�û2��v�`��8�n��tegU[4PiM:�2�]r#�L�ykR��]Rj�C��[�9p�ݨ�faϣQ�᧢��9���%��2�B�� vXX%�X����ۘ����.�|˯_�2s]����C�-� h��ެ�GE)�x��\�@UK^-o �	��%]�󀄉�Ҏ���h��wI���x�G��.�|��gX����p!�(M��N��>�����Ք!|B�f(�9|*�Ȼ1�p`yh��1a����.1w�7	1�T���<���E����ָ�ؔZ�m��=�����j��qp�S�,��2�؆,n�	�#c��6 qs�@��PǷ�tB��2Qk��4�����Sx��~+q���Y�õ���
,���ȹ��6��L�P�m� �vն)>O�����# ��a�ſK؉G����ɜ$�¸�Pb�K�f��u椴���c�0  ��Lw�g@��8�fS��-I���M����:��%y����V2�9�Bt�AIV������\�b��G���"N�Vv��&-2�t�y3�M(K:�{H�x0�0O�
�U�0���8����7�ä�߳�o��J;w,L4�K�L6�݋�A]P�Y"ru ���ϳ��ᶍ���RM�m� -<�d����
��Ċh����Oduo�^�F��Su<vX�M��?��ҷ_\��T�+�#�i���7$�T:��o�3�<lq>�<�XD���9�l�*2�3#Uh�*ʸ��^j*�گ�V�������fô)oa���aC��lF�.����3�C* ��n�q�c/�{��i�22�i�A�%Y
��.�s�Z^�W�
��\D@����!e������^��X��l�U��I#⚅Ro4J�����`�;�Ƞi�ᥱ)&�e� �3{5.�4̑����4�|c!#z�m@@�bf�}����QF��}�xkhȾڋ�~)�ҵ3B��N����Ƙ��'ۢ�zd'�׏�oaFoBP0�R
T:��_�ܿ*l� ��$gR�C����� _phk�dO��*\���L���N�m^h�?�!�w\�+�@�K�R!@�h\������Kֆ��*D��l����P�O�A�Z���2T_>����޾������-0���4��:�tN��h��6m2��@��W�X�>%
`�#,ӻbI
��)��j����1��E���#_�-�P�,,��@���D��)Ԩ���K�f\T'د <1�E��m��������W(�8p|��D$���'��ԑ�|���ꜷ�d�O�i�{�A�Hxވ�tgd����R74��D���}�A��ˎ���*G~�ᔆ���#oj��?K�jD	�O)�HH�_���c�#�7W���a�_��1��F�r%6KC�z�Ue�
rIV+�.��olW����u��p�Ǳ�d@F����sp�X\IfЧi%��WS����/���$�\��3д����L��,1Vү��V/��8��ی�?C���@d86�(�o�5
��Vhԏ̚#���������%��`���([޾ ������]w��!�HqP�02����
K�ndز?��l�`B��C��L/�� .g�L=������:�
�����@�8XI�ٶ9�eC� �{F)�A�%����ߑ��F ��b�~���x�aQȔ��U��@_�b��%�9U���Ҷ���6������jT�Q�?�a���#^{8�3�O�����ף/��D{'Έ͵�y�(+����Gxm5��_si��:%r)��U�[v�4�F���K^����K�P;�'�� ���/WEN�}�	$뇣��B�zh�"�������)7��
(p�5h��b�:�U/����,5�P����Æ`$��-C�}8�>λqjay��'ln��y����� ����c�����ĥ�����֏� ]_U��`��=;��3L<�O�1�9pU�H�d:���'��&7�f��N�R�#�?�5����nO�9{�����`Z���&t��<J#6�u�h�:�_/�߱t�ik�"��3�7IK��՗�B֌���@V���˻?]��_���,&T��Ǫ��F�y�rn@:����n	�d�0+�O��א���E����1.C����2?������7��(�m����H�I�Q.� �}����Gm䖍)�i��s�A3;�o�Ǎa�;]}�{aW�h���/�\*�e�R��^��6k�`ЊK��k��Γ�bX0Yy�g%�����\q�eIW|�� �R��ks�c����{���Ԑ��������z#*�J��\%$��˦��[��i�l��$�E�cR����Y�3Z �A�&�_e��`���K
3%-�L��YF�2H�jf��<I9t�Z}D��b%��$�t����}P(4W�2<d�UWjTF��$�4ϸ��LߕZ/�[ עG�˩!���2�c�{�V@��	�	��ӥ�%��U�NTt�.������TTP����L�����.�'T���v�kO_e�|/�Iw7���ڌ�u���j�\���%%9᮳�Te��x�AK��n���jT��N��KJgX��x��G�λ.���ʽ�x* �5�KD5�O���yJPK�IJ��e, �]]J��P�=���ey18�E5&���~�G�I�'�>.�,��Y��7�fZ���0x��<LbMm#M����k{G�jpu����C����$�,����$q2��:������X�j���n�v�m�w�h9ɳ.�Xҗ�Hy�i(�3��Se&��X��>���k�q�WS�n��<���@�N4�"��e?T����:��7,�n03��Zc�#f 0r��!p�Fmp�%E ��lr韮�+q�k�#y�#��=U�C&E��*b��V,���9Xٜ9���g'w#��9'W�����m�ݍwY����0j~���Kal�S��'��@���QS���pe?�0�3FD��pRm��qo�:
X[Uc�EΆ��,��������B$\ey/�&�.�m��!�1[D�Aq=��[5f��K�"���v��A��y0m�o#N���L�˵���{�r��|W#�ݔ������8,��g���Սy�m������x���Yo�$5Ɇ?�UG;c؎ӆ��<��_���Qt8�Ml�r�������Z���"\^1�JI6��v������w�`��6^E5,
�37�F�ٓ�6�}�g�]�h��b,�>sO*�>���A�[5B
0C�a}��])�T��`����J-�P���9y˔@Ơ]�� �����M���YSL2Z�-]`�H�=������-8"��M�-�I|�1�ȉ�
fɵL�R��D�����I�C̤�`��	��o��T��+�(g��L[q��9��ĘH�$!)�re��q�_��K�k�&���V4���*Z�Z5D�ؠ����CIA<Xcv��0Ύ�oșt/H�������^�d�n�7���8j��C�nqx����&	 �-i�g�(�rT�{�o����Xh���w�]z�u�u"�kn.Ե|�vRe��a�=O��ռ���egA�ΒA�^д$���!=�X@�i��UBb��QgFB�5Ǔ>X̒k�!�n�Me�]W�2�B������_\���BF#��+��{e�Lr��0M��;"�Uˣ(����-�k�K5�Bj7R�J.M�!���ѺHR���%d�i:��"J���c�@��,}3P���Z�=H����aI����� �t���Ȧ��@l�
6h3��N���ae��R�	�O>dߡ�݋����q=������TɀK�L6���dg�.�0Ҳ��%?�.�;�+r�kI˟]$[��:T�At���`�¿�/YK|�N��W&r�7V��d^~��p}9�i�,X���2�,,)rǒ�J��l>�X}K�r�a\��z�=d;$&�K"���2,;Eg1�6B�m����}d�kug$p��޺�7"�)w��8�\�������	6�
�]n	ly����&�Ӱ�n�@h� �����M�{K60��x'��ee�j�E�x����޾f~�j�H#�?08 �a��.�a��<^q>���Ɠ�FU�L�Tt8�yt��!����B5_Tl�3xg�x��Fk5H��M��$ ��,��!�e�τU�M�Q�K@x�[  nO�-J�AdZ���$s#x��'h�#c>����zg�f��!�qCaU�"� Nf�ᐵ��x�{r�/��<���͜Z��quߗk� �`U���J$���N"�k���:��1���p���?q�y/�=��z��k�U#�ov٪�n]F��w�ڄL����~RK��4T��1�r�f�h���^��%�`w܀��Ǻg-_`�U��I�4�L��e����jq��1�?���q:��L��3���Nd���%��%w�|W�}o�����2��f!��ˢCҼ��L|�H+���駡^�{5T%s���
��,�Zڱ\����N��aI��}���K�����û�W!�:��_�b�'WT*�"�	ж�2�UkA�,�{�N"����9�,/���9�`*vq݈�5J7�G�l�Ѭ�¾Q����-�!wu�D��dJ0���m �e%k�&i�
� ^�z�;��x>/����;)9�1Д��*-�����d���"�N�i�Fn�|**��⥿�OxS���wW�(SS����B�ĭ�>n�1m'�⨊��Y��3GͩƠ_�z��Epz�}a�����	�XA�{��2�x�U��[����m"�JY�����{A���U�Ш>o�J)�~p��x��N}� ���D��*��%��7x�7��F��Ѡ��=ow�̢[�yQ��()�ۃ���d2;��:���V^��UH�}��C�ШvU�e��0U=�#����L$����x�E��^���8�E8�C�>�֖F�rxZ�>&ˎ��	bjQ�J	
�T��5E������ǩ��D�~˒���G+M����|NY	�=�Z͟�4����6ة�:╰^���җ���3~k�5𹻗��#w���
g9L�����P㭟d��;=�Q�ޕ�Ê�9��˕|3rΗmc�x�9�U����-���̘�z~02����l�	��W��r&G���Z.����GX�j�t-��2u����Wp9�o��`�z��)��D�����O�(F2rPټ?���C���y6 �_���;�v�uO�6s]}�i�C=�^(M���w��b��-!���&.;2�S���N)��?�Y'���[�=-�1�p7��A��з�$�)?C4ޠO2}9��(,��|���Q�8QH��a*_u�9�gc?�۬�WX���L�4	�+BL^�f���K�Omٛ'[&����4%��
~sk� ��3�b�8k%���YA�fL�9���3r�h���ۡC��3�s���wѭރ�9�����!4�sD�"w6z�$V���Oc�[�K�w��ٖ"Z���,*����!�|8��K�k���Y����=X*�v"=�7�� ��>�A�T���a��
^�����rAn�!wY�tN���������dʚ�Ҧs�G�� M�Wl";����ǀ�U�o�� �g�
!,W�Q&�R%�4y�j(���0%a*Qe��g)LXhV��)���i��v�^q���}o�l]�IB�]1�@YCy��hb���r��R����u]I,�J]�(����U�̰�V�J��$Q�~�~`<d�PM�V����p!�_���?݀a��&&��+ro�[R�H�6��j��O+F�c�Ͻ�������=�����$
q��D0�W���&�>ͩ�] ������I�S�K<>CD|L]3Ô�?~�����#�k�#~�O������2QI>h lg�s�QF��r���Hn��)�N\�bb��@�?����R6~�׃/q1��*��`��}�U F��a��ʵ����PqE�џ���e��U�*ءh$��Ϙ$浒9^��������F������Sg�*x���mEi�{DsZ^�V���)��|ڲ2��xu�E��I��x=�hKo��s����	�7�h�<�'a�pӅEKrA��T�Ur#��hƟZE��R�t��"�E�^/Htc;�b��q�d3ϰY����jցrY/���(����>/HX�[	�_�L��W�/�ח�� l����V��/�G�Q�}ָ��K�lx�I��ț�#��>��hi?�I\:ُ��̱�1B\�`Ȕ�¿!������n�����)��N~����|O����W&��|pB �'%<��Dp��,��w�� 6���AV'�β�.e^"�eʍ��7W'b�M�9��-�c�?�,�0o����:i��k�V��³b�|�=aj��n�6���b��}��/8��^ŶD�3l�z��:�z��� >� �#������E���ը��E��/�����������'�IkG.���Q��_/��љ޵
�VrF��4��i���b��-��bɚ�c��U��3=����b}ux��z��hm��-ɹAt��Su��1T��Z.�oȩ��`����F��{��r��4��~��$.��B镻����Q�m�������R{0|�`�iP)H���'ղ�}?@��)25��(:❩�ﭽ�V�G��6���s�y1Q���bh6��R/���� 
���Pꠔ��Y�1]��k����!w�3T�Q�N%�0mS��)�:���3C�~�LN
��r4����\FZ4�kç:�g�,�rkX��C���(_"�k��3�R��b8rV
+� �2g�(��r%$`Xt�F?���4��s$K��,�����D�9Q�Q�S�3�J��1�⁒�_�K��y���ҙ�0z��6�7茎u=�艬\n1+�?s�H2L1�/�ura��jF�4�w�E1������V�=S4�`Y�e���¾Ck_��]"����J��*^-h�0C��TK��c7�X��s�����L(7z�6�E\94$�f�b �k��e�g7j0���:vJ��u^2�\!6�=MrC\���s�F����� ţ^���H��,���E�p�<\��/]Gr�}��Z��f�\=Qb"��9,�3���5谎c'����e� �6:��?��C�����*�h��o�\�akg��gT�bD2H�ޫ��|t��g}m�J�;M�m���#V�{��,��K�R�t���_h�E����/R={�a�e�d���]u�EpӬ��tu`�?M��H�����Ē���e��k+TW3$,�ӆӡ#���O*�E�y���5�N�Z{�)(��y3kީ��?�KT�(��UK%���?y����0�n�#5����S��ۿ�&z��X�킃>㯈V�����E�|?�K�M39����=�������Sw%N�����1O�������o�ѧ��N��U*���b;�`:]�*9�E��-�XUW��:��"���Z8�Y��4�!�+���]}*��1A��H��&��_i���h1)���Kd) UG��K��,��F���O��E�N(�B�`�aXif�Ga����)uM ���h�6c��-�z	e8���1x�	x���V�S�o�"��`��N?�z�|��nruA��[��.}d��k �Y[-csu����e�YS}���'-BM�PL\��Vk�u�#�����a�ț���}N	m+'��U� �!ȟ����m�j�;�-��j�MI˞��9�j���=2��-���	\�[�xN�ny�ꅦ�{�|bg����ّ�\P��n���H\?�ڼ>����<hQ� �ٛ��T�n֎��O�8�5��ٰQ
v�޹���u��=��eQe�1=S@X�h�TJ����>��JH��q%���\�b�yne��X�A�SA�'>*����qH)���z����s��� ��,D�����ݔ��e:��*ri7-���\��ۙɴ5�Ȣ��]�,6��x	����O^�A[�*_	��M�ȣ��#�^ ?�'����Acח�q7UY��ݡ�3C�~��pD��@,��>?�[�,0��B(%DY��j#-�93���'��Hz6. @�~P��qNk�1��b�(��K�R�r��KA��MiR�S��P5���˽���o����U�:;%�;�,]E�	�g"��xG7>�H5�
K�x��S����S��3}itp?ŝ��H�oP 	4��-ћ�%���ʃT�ۡ�{G�/��PE�Q���p3j�6�v���7�5�TX�?ad|�1 Xw�!��AR�p�s?Wh�|L��[����]�X%֧����q{d���x�V4l�3_�^Cи~+�f��Y���4A�Gs'�L�V�9�>!�N��A��i�˙|`47ʒA�G9UU�l6$4"�ˈ�В���&/�L�uⱺ��IZ@�`AC
���O�϶�ç��� ��D�lS\3�}S���qםЂ7��`'�l�4,��bR>�ևc���5.Z#Ȅ?	��e�oLZR��ʟ���$� ��W��!�R'��ʅQ��4�W�I��b�ң"��c��x�j�JXd&�f��F�
�N����\Y�q6>; ���,h�<]�0ӷ�i_��!���qHrćo�'i����V�6����n to;J\����Ud����m��5a6���F��E
z�L����/�L%M:m�;�K����� �Z�شܢ!4B
&�3�}~�O#��z���{UL��������_�rK�b<s��L���s���I��%A�\��%�TE]��S؂�d��_��2�I�j,9���n�0���7��Uhd���3�����0��2����	DP0c�?15Q�X�k+x�̖��n~���KBV� 7�����	�����#]�F�t�����r�ؠ ��/]�WsζAD�8�E�����!�b���">}�D����<V�@�I�zM$��I�v������yy����||���j��,��~߃��G*<P3M�"F�SQ��>B�e>�����з|�dE��n��e
�'��o�8�T�n�_%�"���a$/6�TUfya`L�R来�����qB�vð�io���9x�a�	��g
� �)2��T�eo� �&�����1���2�8��?�Q��TwQ��U��娻��_q\lvܴX��]6��ve�}���_0�#�t��e.hM�]�S��*`���a�g��+����/J����ZTA�`��m�=l��'�q��n$K&i2��Hf6���9xl^aﭽ־_�n���|uC�/QE�cV2oE�r  }8�p��>;�-.4�M��K�"v����ڗi{�h�Z����!��i���8�U­�����g�#���=�N
�]4��N��V�S)��7���Ɓd���Jj�Ce���J#��oih�_K}��xd~y��3f�����V�����W��C�^��F��Ё��6��a �]�P�v,8c�Y:����Ӎ���\�����i�l�C����j�VA�C�n�L&�D�bxߟ ��Х�ɨ(��q;A����������Z�6�Jݏ6,��J܃>�ZJ�>��%�<��ްN1� �7�xm}"�ˤP���n*���A�V���ә��͏�BF��S����5���p���Md�}�/)z�6�|�`�*�8��qբ�����)�#ij�o�e�A��HN���z!<u{�M��X1�8XS����ќ���˲��U�?�|w����.hk%�F�{���.W��n�e�SI�I�Z���Q��Z���0����ُ�� ��4U�kgBi�W��H�Vg��F��6m��K+�;c�ڍ��&`�d�,x�M\Qm�p7���X.H+�`�����|o�(x-��σހ�7������5`�Z�!��IED�2Q��<z5���'.7�q�T���p��_�{Uk
�&(�(|�;���#��O���y�1om�9Zy��#F]ad��Z=�3��6��S1��NB:t��&���e>&(��&�j�@q)T��얲v`�X|%�j��D�!Bk��#����W��4%�UQ��۪�2
�s��̾_�`�Sѡ�
jqN~wN֮�����2$�����b�kǲY���Y���r�A¢���f��NO�П��ޙgSn�N�g"���5��N�=�	�릹�����]�������q�����* �fZp�J�(��;�Uv䨻8&
v�`��(��}�GD���;o�F����-Z&�F1�B������ZqKМ�{&�$�*L'��[z�^���Q��A) �	_&cu��$���ϊ�<����$�Z�'p�v�6#�WsP��LA��}�q��<x[��٬��t�GJ�h-��VT0��(��Xa8� c�$��I�"�n�,���6�ۆ��mi1�S�5�-IR���~���P�opx�
�(`Jh�?�ܹ���}�H�ə��/�0�y�������N]}Fu�v|�a5\bh���,�Q;tz�-3�������H����s1��,l�����
��@���\dNB.��^���x\Zj<|���&�]��/s]7�	�<FX��|�Odܖ�m���o"ɭ�����+(���`"�V/_�����?�N��s����� �Q���H��C���l1�D<��rf3�p`S��ι?-���J,��T_��C�Z��K$p�\���;�J#[�J�'��4�m��E`r�������ʅ�
�^��d�:�b�h:6���x5��)�)�~x��G��d����H�q��U��n�3G2��mm;��T�EG'>D�F�D��R��?mPd��#1>(�<���h��̿��[����}�*27V���\��k~}j]�7d3��4M'�?1ݭ��ɮ���X�C3���%J
F�qi�l�����?��T+�]ԉ�[5렳!�����dC߭�:�6��t�`�._��*[w��e�R@�B�щ��KT��)q����%�o��Aic��b8�� o�lE�}&<Q���� �ۿ]�x�Pc��uwD�Ќ+���W��-"�TJ����.8��U;e����?jw���{��F��X�u�Rd��[<�q���Gj�n�<q�P2Pe�5�"���/��ґ���*��A�l��5��)8�תN��=����M���L��߰��q\c�X2�*�|��l��d�t�;r��c	ךr�1G�)�Z�`����$Mu�ؾ�
i_�r�
�,�Vh��C�{����+csS�[	��5�OP[��)���Vc��M}D�'�-��|��G�����ㄖ�>�:���W���c��	�\I\sT���������Ӡ�ݗuS�-�^N�#��r\L0����� ��_ԍH	�W_��\u- }�">'� ����=5�����B��ԊۀYN�t�|
��M��I��T��+!hɦ�����F��U�U�C�_���( ѡ�≺��|v�-��[����������w$��e�l^�b'�a`j��#/�M�%5G�Q��g1	��Q����{\0� _�f��i�\�x��\4�����yb��b]{ǧ�iW�S��Qb;U��|���e����u����djK�:��3�͙,�	���˗:��|!���z?�����԰�B�!,j6F�o/<�v���G� �5G��ƸE.=uUY�mi���g�y*�j�����?;ޣ�KQ�~�"�*�Q�m�C҇xr�5+캵�	��@���kS�A��Y���^��ӕX��PJ�H�Rw����?D]��A�2@��"���4-}���v> ��v��7��X�MR��'Ӛ���$ݽ�{Bޫ���$�1q�z
더Z��d3�����U���}����y�VIҗ��C���i�\k,/�����O��-��
$��j��p/�ם�~� �?A���O����lShb ��=�2�N`w�Վ�*��ِY;��`e��bK2M�rK;�}�}��Ia�<���򞌄s�p��7�o�yũ�/�*@��������X�����l��穓wdUm8th��rޚr,��%C�D+/�*���3K}�{��C��!j�e�Y[@�
��)r��}u���z���2�k�����I����*��e�C���>��L�J�ӯ̋��Bm�<G>��v�n��Djֆ��-�>���	2
d�������6ZÙ�J���=�"��ٿ�خ/

�ˢ���˥璟�� �p����M�"����A�T���#*Ru�t�����`�6t~��ěc(hq���b1��uq���>r�>mު�����D}�Tɚ�[꾸�4C%3$T�s/쏇zջ�$E�0���%�f���e�yjE�4�Z�<n��wl�;�ܨ`��2��[_T5��U@����d�[�B�JC�@{�45v�������׈���K����+������7�sp	e2��>(��9�Q��F-'��y��/pʚ��V��I��4����.㥺?��zQ�Z�*��U���-�A�Oe`}l� ��x��d	�=�d�;�5l�F���78ۄ���|q}������r-֘8A7���0���O�6iۋ�EM6YW
�0"�Υ���>8��0�V�7~ۭ�s8����Y���}}�F'��7u�a�-��s���������@�:ĚaOy����7t�\�i��m�KG�U�g����U��(� D�B��d�Rc����F`�q����������X]Q�Z�B�v�'�Nb����|�D,�r�
!�>ݐ�hU��x��/Fg��)J��ZT��MZf�]�ĻSQC�{��B���F��W
�+r��]�\|�֑9T���i��'�l�xC� �OK�>��Ⱥ�B�;�� �1� l��EC���*�B&J_R:�FuGUD�J^eH�������=?��?�{�;�F���Ǎ�n��_��=��Q$�jI��D!o&�G�z>1�����j�%�A���5�1O�#,���j
׎�!�l��9/,����1P����Avq�. ����g�@J>R+�X���N�gFzd҅�%\%(�*��\���T�_ؽG�r]�Vk��M���Ā�)|��t�E)b��&�'���p�P�Jܓw�����n��+�N�H� l(�.9F�0�[#��g����̫*�45Ώ����x����o�N�v�u����ą ���� �+4��3��i�
����|F;�y��ت��'�P뻉�d��@*a�7�$J�r��e��W��KgŐ�DR�<�E��D\�������e�,4���3��x�o�g� *���|�y�o	sϑQ#%/[.H&8i/W���-��+Xq� ��g
y�9 thI�I��UZ�ȩ�~���QU�b#9c�t7LQdj��7�+�Vs��}����4�{_itE���?��/�疀�amґ��0o�r��ϤS�9���	p��q��"��1����)�$8ṩ�햎�j~hju~����q�zc�>}q��D53ۚ�r ��8":��d�Gs��"Ed���(܋L���ȍ��SY��l5}{O���^��0@-4�|!�žu�A?��e*"xWW�he�gĘ�9�����0�Y"�=˾T��T#X�3��qly$�m��!�O�����,��s����CJ�f���!& ��.��6�K��= ��F���������n�6�+�	���|=w�@�4Qol�V��0�ٺCݦ���+8���8��ٹKj��T��]�>ߵ g��f���Q9₳m�dx�C/��h�{�$A�$�]S�ٻX�SS���8�9����K�_����n��k'�Ӿi"�l����p�
�En[�Zoܐq	�<�'XpUnF,����۟-���,P����^q�ʚ/��6�`_ϛk�?�x��z��"Q{\���ש����F<㠿����h%bH���r��OF $��K�]�����Y��K�T��JUJ�c���[&��y�8
�y2,���(g�BK$�2�;ɹ^�� ?��?\�JV�ڌ�ț�Kq��R[���+����� $ˡϺ������i�T@��b����>��V�\��L0wVDܢR?D���RrZE�g%�k��T�h��Yo,�'�kj�t��4t�j�(/0���es���2������%�I%LmW�Y������'�F�~���X	`�x��Unni��� �����p�����un�UM�T7r�p�i� �V�Pp�	q�%�ԝ�i=R��U�G�I��iK^�RV ��SR���JV����	wn _+ǒ��c�*�U�ٵEm��F����"i?ba�s�_�.��L�>��l��M9��$j����!D�H�_4	�+`�u���d�C����J���u���{Ad��e�ڢa�͘��	s�N`����p���2̒Y�%�����FjC�P�Ն���K��3:��	���Q���Ũ���Z��Wb/���u�5@�G�d��m�֦Z�?q]q���A�Ew�CkP�����EJ���^��vU��4� �-tCO���'�9�V�,��-ʛ��8+��`l�����22-w��c@�<��e���m�~�&-������K�L�@�,�����D;,�!��6�g��/SF/O��$���~vE���Z�I�egw���r�ia�����6"�%Op@a�<��8�r���u���&~ a_8�Yℾ�%�-��n�6�����&I��)�/�����kE�<���,����г���0��]8]�B��x�qs���\����A�h3����['�#�ϫߡ07"�~�7��2���#�-9�f��՚�n<��������J�]P�c����*	ëm�|}&�<3y?�# ��:Km���!n�"��L������yk��pcg�ǔ�K��ԟu���zς�wP&���aS�Ayȴ�q��񿃈Q�w*czY�`�s�-�-j)ja�����`�f�1��&L���ܥ��;s�L� @��B��x�ydĔN�ލRD���o��ߜM�u��e�!�H�2��z�I*44B�aq���t���T��>�,�b�<�!��mlAL���"��_۰4����6J���	pbH������OxQ��xS=Jg���5�&~�%�5w�\W|��q?�bDwޭۈ�IPp�>�Kw��"�/��Ia�E�7��.h�W���Z�����jMG�мطb��h�%]]O6�LB����{��77�)�8q���kR=��#��7��#\���Z�=h�]Rb��@�v��:�=�J"�I�����U�lQ!�V�����$C(X[Hz���y�p�,� 6E#��Q���|�������sMX��U74L���m��B�o�G�Vc�::���R>�b�,�=0��~	_�s��[C�Ǥr}83i���[�$"6	2�/?nSꓟb+#a��&Ʋ�{�$�)�4U����s�m��2�!��D��I=x!H�Ģz+�l}@qB���|$��?�T��|X�L�ް�؜5�g�@�u�}z�r��Cm(����*շ���hT"u�	�M9�ߣox����G������ �$�-�E?fD�q�=_q9C��A�h���X�=� ���C���Aȗ �T���R���0yu���f#��fZ��׍q�t1��8���E��A`~U���z�?̩����"y�S�vɠ]�͖uэ<������������YnUY�|�|c������]�T���h��@5��.��%[��+{M*G��h9_��,�YM]�?�U!���g��wG���ID�~��_]u�L	�L*��7�	�-�HM��#��q����4��I�m����gt Y6S�}p��k���bx �3�m9�q��<���"?s�˟ �uF:��4ԭ�b+*�B��~T�2���r��8���{�����N�x�'���P;NM�x\|tuz�D	�x�7��S-u�^8����ܘ R�m�qj�m9�t�$�G��pi�ot7�hb���*��N�Z]��A���Noh�2A��� T\����c�&���q�<e?�$!9_C���k�=u)���=,�Ib�h{�.4������k��� �ϙ�6m�Cs��)#W����qt`�V��/�	&S�Y#i��R����L�v0-��yv�5.��u��'ذy�"�S��3����ܸ�c@�'�&�68�c���B�f(�4�ayrW$@ K����W����x��<��-�.B���K�z8�]���M�ί���)�$*�-{�_�n#�x����3/pW�'�Me��E4|_mL�(t%f�-�Q�V��S��ê5C�B��4mN٪MY�p��up�v���/���A�<��ǈ�3"�_��ħ��I���parLw|�HHC���t�)�Y�bf��������w6��o 
S�%E!�H�RDs��s�y�3\녺	�/��'���f��O�f�n`���'�l��ޔ3tgYt'�����#&7���/Sق`yCO��P\
!,�K�|m�de������%������5M/tu麛�n���d��p�R׈z�X@[�k������aa���l���"J�~�S{�7A�zgM=X;asǷ���0��kN<2�%��B��f"�Wa��d�h�r��)�1H_p�Byp��A=D\��C��a�R�6�^��Y� �+��ل*�������@���~�`��Jܷ���@4���cqπ#l�Aj� +�x�iŔi��>Z�
?=C�Ҳ�J@���D�zM�̬M�.*���dK>����9�d	xće㕊���6ZP|Y*�~Z���:�>�� ��n+�7�}�Y>�涱�{� E��v<j�����@~�l�f���񻟅��v&PDhh�+�HD�ע�8��N�E�%������-�k� '�e?�fC��1�,����}4���K���湷�q���B�����eң�z0{0�'��>�_���V� �,(�3����:Ug�3��Z���S]�Qu#���9�v'mN�v���*�3S�%�=_'�m9�팦���.V�u�vϞ�T=5K�wR`��r�ޓ��IJ���q�����Ï�α�4�H�V/|7w�Qn����[���5pܚ�!�Z
��"x�		����;�7��T#��E�'I'H<5��ߕ{ )偨;י����;����G�A-̗e�%�ҜPf�!-���sZ�rN�V_֜����;%��GX���tZ�Ƚ�O�Y|kՐ�IU�A�̻����iպr���W�����&I=�)U1�'�-���� a�P��O��������FF�aL�|�m��iD��M1V�q�Z�I8;��D���;���N����p2���ztNX�ӨVV�$Bn��������Zh3�#�$E+�ʵ���A�qZ�4.~�Mk�1=Q)Q4�����&�I/����Ǣ�5�H�}t.T0���>���S��`@i��/��̳�ݽ��c&Br�6�6��-�Hz�9��uN;o��A~�DNY�ݦn�`�d�:Q����K�Va��E��lxVB8���JMc?���T��Ё���q�D���.�R�g�,�~5�����]�r��h�J���"{cy?�w����n�m����[?򀓉~��piJ��%N�u�$�?�:���B�r	�ZE������r�3�Κ�F�+(�Ww�t�/2�i m���G+�_/��~$eRc&[�:^�u���y����#I	���0�wũ��˻zy�����}Aw�sGܽ+,���3�T�F'|�AQ��	���C��;����({`��#��&p�p�Y��R����%���aóbj|��ګ�%>ugl�#+��eV�af�vX_�/I��(�5��?Tδ��e���y��q9�f֖wb7��
�2"��4��G�l����H�iP����Q��	gz�tx8/��J0�?څ�Kfm4*�8��H8����x$o�Lh�$�8~���P���_Md���75��09cd�3�]U����u�>���Vʿ97��y\�v����4��]��Y���O���F����aU����ef�XT�`�6�����v���m9�dpfp��RJl-b��,����Ƭ�~���]Uwɝ�L �
�6�����Ō KF����C=�,�a)���Z��Z ^5c�Hq��ǹ�U�l�g�Ȱ����
��Oe�h�K*;��^X�K� h,8semc�=p�)�!�Xg����ø��22Dɿ�p�8�������14�Z���4e� �ϨT��f]m-���������3-�)��S�-	�Im����o�g��c㘡�;�/#Ů��ܶ[]�=�\$���V���T
������h9�{��.�Kdf�R���)��c®gE�|�KP
ltz�`�x��C4�yc�\{��ey�Y~���1N�<Ӑ�U����x
T!��%�<�!����ɕ�� Rq�Y
��u�4'6��G���θ��*�):�@<�ҩ�.}�+������v��x�c �Ja�R����|�_۱@�t��{#�uܴ�� b�w,�7���opqr��_�<=��wH�>x �o�g	,�n�C��כ]�wZ�����0録��)��^��rb���Wɵ,����O�~�z�甏���V�?'BE���$ېhj�m��ph4���T���*��e�Qr��G_=?���`��n��l�����Wfmrl#\�y�)��m��K�
��.�F��Lr=w�)�Gl����l����iSS9���]���0�\8;	P���Қ��*⫱>�K��;�0���,���f����%>�;v*^�ﱈ5�-I�5�f�uׅq�H^GlD�ɩ��%�w"���� ��~�%\�'s>���O��Zk���Yn�g�h��'e� �ݎ1�Bw(ɸz�e2�墚��UO��F9-�۝m�����}@����V*I��O� ǂ���;�\�&v�C�9R�;t���8�`��f��Y�xc(��(�`
'�.��j�_�������Oej(����7" jF{��)"o�@%�aZV������P��g��D1:8O��d��ӵ�����ў���a��u�����H��`�����!�Ґ�tŹd���R��a����2W���ϛ@������zL�?�X�c>�"������\h�T���q�߃���u�ܑ�~}�Y�B���&���5���hG���?�'ˣ� 'Ba�Bq5'��	͟o/o�5�`-JZy��@q�mH����^`��xsQ�?]Ѡ0�l �Yx*Ճ��b+IY!]֐�U���P�P�I�EѸ���/����J3^�X�
�8B�*�$Hkb�ͱZ��D��Q�X�Í�;]������s@����Ld��Er6x8�[K=y��̯�u�k�^E��jL��v�l:U@��&o��?%�I��P C�v_�������g0�z��b��m�j��1�.��l���Ӣ喖e ��|�%/Me���g�8G���9q���hKC���I��υ�N!���./4wd�X8��U��a摦tP����Lկ�#9B��1\b�����ĥ$���~e۳���Q�՘�m[vS��kkV-,EO����e<��j��(*�-o�=]2�5������s�/,�(=�'Q&V���|�24���-��N�2��a_���N%I pĤ���G*~W�cv��	^_X�n��i�ֈ&�$-�I�`�prjl>�z�DQ��ƾ��Y�)]��]�C�DY�����ev��c�G�џ��N���:D�_���=L 9�p	3��7���������7�T�r9�^]:�'��S�-�98���-�a�h��Np�8_K`I�s�y���׈��[!��ı�	̎: ���t�&��!A�r�̓��Q�/Gz��`.��v���S^P��4	�P w�[~��H�i"�<��j���+��%8�9cyB���fa�-Z:&Q�j&���ey�(��|2���e�>��܎/F9S�;�1�MX���w;V���D��T����$�.C]:��<_(�����&�vm�5���l����9�8��G�2zr�z�Y@o+Z�r�߷�9�7��f��o��R`�W������!���@pI��*O��;�PpLT{&�6	��r�/b:vK=n���O��t��)��B���4� +f2#X<�a��7�(Wʾ��Dr�JUMVu�|]��x �Uo���*vcv�#mlTO8;Bc*G�܍�_�ա�פ��vMl�G�9t����I�sq˴~<N�'j���I�<V�e��H=g���Ȁ�R<5�m�2���U�G,{�?�����]��du=��MhS�[`��L.�Ū�q��� +g��i>��w&�(5�tY�A�n3�C�vAu�Қ*K�IW$�z���}��/~p�wI:���,2����f����b�C�$Q�YC!H+��\��N���%�p�g�(���E�77�
�B&��gG�q8FW�ۮ�����rBM0t;�a�Scazh�o�R���E7�G6��Ͳ�?yv雼�Tte�*F$�BWpd��+)G ��p.#/��(��^S{��F�aXA��$ϖ�Ϙ��Ԩtr��l�,�|��D]8�X@v<�'l��r���̳�,\B/�/��u������[H�3��g������|[c�#y�D��J����UJo瞿�ßw������挖q���eb\0�A��Y��V��{�e]16U��S��yH�)�J��3���`l���n��Q'�����/Srp�B���(-E@+�i�37储���3?+y���T��o��?U�WX=��~1�J{�4��o�:�5b�����m�K��K2�ݿ��`���i��N@M�.<�3���2V� B��,
�A<N!��|�ӭ\�\H�� ��#�/�@��Mܤ�:�x��7t^�	S$�F��Ԯ6�2!�?�˙Ю$�0���躙�+&�8�a穈�����NWx%�s��k�1b��nyr��^@�mǠ3Ux����|u2_�Qa�5�x��f����L�!�)��7K�)7[EK2�/�6C��rl~�h��A���}� u>����m��D@�F��H��5��K �fV�XEO&ކ����ً����?��O��b�mTKя�9����!L(��{�\�%�$�K�>?�� ���V�Pa4A����SQ�g,����C�]Vjbp�l�߶s`����v�����ɯh�[�+���Ԩ����˗S�S�A��8�j��q���-lO��G�oW���u1*�^��޾M)��G��ąQO�ѹNUFѠ�)���������J��R�ܰ����K��k�:�ױ]=�l����1��(� �x��V!��}��"���K�8�xvD�Řx�A�jR�K	��i�G��2#�u)t�7��2��3i/<ǿ�	7M#�h��`�{,QL�8?�%r&4�#��~R�oQMM�W�<����ݵ���{L��,��8UwV��p�%��� ����dт����0�� i���ǁ@�z@�.](,�v��]��K��т��5oܨ��+9��9NR�)Ģ��i�=���DsbOŝ�F�C/�m��2,�k� �J�c4}����tA��q�?B�ѳ���k�>�0��In%�
|�����Ȇ!�Bd�D���5̞4P��æ��[9�,·���$��I!"�]��s�N@��O.�%�H{հ�;���9�|veϤT�X�ࠬF�GW�6���U�A�-�-��U��d�V������;S$#S.���k��hH����4��)?b�+��=�3��m9�v�.�>`��`�yu7�Q�U<"��!R\��#d��R�e-CC�'^������nw��R��R&���M"If��J�����6��M|?ӂ��u�y~Ɔ�^	��1A�Ѹ�U�eX}d�hӡ:��@�G4��K�1�#'a~7e�[~G�RJ
}�~rtx�?�_.�n�w�;��[;�scc2@
��<��@���B���H��n4��&g�+�~�m�]%�⍘ �����-6*�m�6�Nn�N�5;s�\=V;�6s�,�E��V��n���� ӅD�w9:�3��|�g Gf��#c3������$�1r�4��8)�b�8KeƷ��NE��e}h�T�����I&xmt9�7IK��IH���i�4QZ��*���PrF��븿���DB����Mw�X9�aj�x�H�ɞh��<����3�H�[L&��iҌ��Y��.�k�7��TY����M��]��zצ�?;7{��{����{��$�ǜ�:�`���z���T�^A�o�^�6��7),D��ۅ�JH��z��ѫ[ ���DG�r5�A3���5�t.�Q3�^�;����Z�L
��6����`�EBU	���Gƅ���
\�'���v�X�.��tv`���_���5�0��t�.$hh��9�����r�-�uZԿ�]���������e��A�l=}0�rf��R�v��}G
�1�{�;]��4��V/-�^2��+�<��8	Be!����P�q������⚠��ff'ڥ��[�/�1j��x��7�`�8 E�$�
Ŕ���}��t`co3����~�@��v
ex�Q	�N?�>�����$|�Oٵ�m��gt�h�r�K��V"щ�ܱP����*�4�L�2�v��|.�j_��g������H���ug=�I�����t���D��i�l���\�=r����4:�CLiQ8�����C��3��#����eM�zhk� ˭)w�w���j~�!�)�&kc$�lw~�s�H��>:�� %�}�u<Y�~=��L<��!�g�ΦUw�udc.��B�W��b����1��6��}T�X��!��T[�1h���b�/ǧ��Q��L��'�p����o���ߤb�,f���ӕ��ʕ�$�����8�Qn_ArN�OG�(8����.=��~��4�{��f<8_<�i�9JOr�<iI7�$��⧿�;��97��mh3��G�x�_.j�V���O;�i�w[���^�I}�Q�+�l��L��с�)�筕t��qӅf���ٓ
@��V�f�Р��� �~���vR�0��aw��#��F'�Ud{�g�O�vi0?���ͷ_�����<^X�򜟘s�G��cp�2 wL��F���m=q���r��E\�-t�ZR7M���ʵZ��9(Hh&��G2n�BNfI�:�X5)В\�\�91��*�Z��U�F+��q!�4�I�!t8�B\��.����<�2'h�?��p��3����+��m|KM ����K�1Nɛ��ձ�Q�C0�
��&FV%Q��ꮰ0#0�)�/�ԁ��e�;?�K�ۯ�4��,	X@�\�����\�����;�E����j_V�	ǂ���.;�����c�^������,6�Ս���u� M����f��)Kt�0������w~�*��c�Q����l�t��E=W��FR_~�
�I��<�N�ڂĚU�V�#��H��@̀��C�}{�*j�"��q�5rn@���X�X��H��~$��R/�s�����В�W�^����	.x�1��̱�C��K񼴖l]�.L���)�����aX��ֿ9-$΍���gõ����ؙ6�b�)s,+�W
oV�۫I��iN^�S�H�3_;j�.}�)����B��xNQ��\��+���
K���_ۢ�,����d'Pl�;�+���"=9����g��6i!����06�.n(���%�<�k
Q�h�[��iy�5W�:�P��Ѩؿ̤ͨo��evʧ�>)�����>MA��_�$6bY��3!����J
+����D輴z����eI��!|��g�e��C�"M��nEzkp�b:��,�[�W����������ٻR��83��m��E}���؏˅-��89�Cz�n�oCp��D�UKaA�<��I�+��\x�Ύ��8���	%e'��܂�ucn���cT*4Rp��hl�"���s៷\ �O�A�z�s,�x���Tu�:h�q��]�|K�M�D;������S}5�š�g�E9}����a�n;uNbuK�U+�f{X'���݅�O�zM�d����aF�	���mcOܥs`�L�x 5��N4ܼx-�� S� ���2U"p���Q�����q��e]9��b�j����D�Y�i�KC����I�(�Q#�7e-3N��$�.	@��������DIO�n_'��d�˒,)�A�lw�����ᒟ*�VKYY�չ�2|�b�W�|���	��I&���&��䆰7�9��oh
_f ����t�&�^��m2�Z$��0n
c;�_a2�VQ"�Um[���q�vMq�?�㨡���(l�4��m5�z"�L����2�[7��Z�[�����x<^,����w��F��D�oj)��y�"��-h�oAj�v�0�3���\�룖�!f�\ss�M^�Z�9��?��$EF2�-�*�*s-�\n	�`�;`7�uG;lWˑ��q#����4+6��N�$3M�����%Q���-}W�/����[��$��d��ЊW��\��1H��R���G'�O-nV�˔d���]t��\�HN��;��:d
h_<�&��HG�G�������W
�m��w�t#tgO��i��/�
�n�w��
�]��Z����A��ϧfʺ��-����3ÊB#��S}���}Y��S��g8��_[�4��4�������0��4Q�[��>E�/��G/�{.`y  m �������s�J�;�ݩ��Mܣ�����y�X�����V���?�~�4h�_�֭;v��H��4��%j9���{q2���:������_�-Gj+�1�V���9BD8�
�L�`���	u5$(��zR~s�]�;/�ʹ4Q�����Ԓ
�}G�M@������Z�OCO���1*9F��y8����=�iJ�r�@zlF������?Z�7�f
��p�VM,�b�;9��}��ӟ&�����J�yd�����p���y��.�B4�E/7��Wg�X3h��RI����k>fV���OԖ�`tFv�:{Or��Gg>zlU,m��Y���`�W,� 1jQ��˧f2�VV���ͼ�c �f01>�@ҳ������C\9�Wf�y�EB���/@[�^[B!��gN�!˭���i����{����uW:�NȶRV9u����)��mU��Wg��2���h���}�/qp����~������q�T���j��=�b��\#�����Fr�L?��ZTp	(8��|%4�+^���+��#��U]Xo���Pq`c�ׯ�q�^�l����|D$g]�k�L�4eJb�O!Y՜t� yK)��͓��y�c��U�_���h�(�i�R���8���G?kIbU���N������q6�8�Gvu��Q�"�Q���f�̐�^����П��`h;g4g"�2)�c�7�#%���#�,%n�6��M�#?Z��O�nf3���{�|�q�-L���a��s�-@:�c�E$���A8���Ed�y2)
���v����^z��Nc���E�y¨�!&��$ް˾������u�`�v=�rE��|�b+�K��^
�v:��O��� 5Í�k_j�t����� ��>�����vL���Fc Yi����(�2���~�k̓ɗfoH�5�4B����ԥ�B&�������ͪ�>,ֽ����Z�:;1�J�O�}�{���'�픆����vP8�y��!H�j�rvP��agJ �|v���1�^(�C�#kQ8�����Y����r����pB����of�\O��ZA��I�7T��g�n���eP*�,Ξ��Ǔ���"�_��dY��Z�sz������j<�O��v��F��;�ζw��P�G�c� h���P��<���ȡSb �s}������<i���@��yR9����Kr��Åk%���P+4̛
���b�Dv$����xP�JT���,P��q��o�rN���(%��$'�VGpU����X������U
Ggb��J�
�D�=�w40����!On�O���H�����X0@f�\���aa��T&��KR6�#�H�J=&��D�k�]�HP��9�:��Jי4f6�eA0`��
�i�A�?.��� �7�+*�����o�1~F�P{�!�)rqÝ߅���<D���T3�z��q��Fa�Wq/��d��8�J��y�bh*;Z�g2v�Z�2��U�AZ��n���l�0���-Qm-Qb?�K���z�����C_by~G[�t\a4h`� H�h�����T��䝴>����N!l
d�\`6{0N�-Q���b���3nd`߱��r��V'�e��|�#��Pj��׹�T>z��Փ%�����}�q� �5m���$���j�)�`C�~���u=��0�Yv�Ο�ǂV�7[aʱ>�~��l�A��z7��]�'�?�1q�XS�l��GҊ��$Z�]�iWmh�YG3��u�cH�n
#�Ysg����3P� ���!�%s��ͻ�L�l�S�<O�:�4���9!��	���2w��l��Ӊ�2�#�1��*4�K����o걕<�1'h�7L�~9�O�����B��'����<i����y���vh��x@Pm��Y�6d~��W���LH}c�����I'�7Z��R���/�n�]�T��pp�2��@<�YlS^�_��5 ���z�J3e��W{(�uX����JT�=ɍ�0��d���!��Z*7~.ҭ	݃]�(&&�7^I�V"Z@�@,�Mb��
&�c�(~ఔ����m�3|��r���9j�%��-��}�6J��F�PR��0�"(�P��,r �t�|���,��V�%Q��=}rJ�T��yJz�{�ʪ_P�����+�]_��x�_V��w���4�b�4���ș*�(d�_~�Ta4U[��vt��ތj���R��w��*��f*��r�h�'�te���+d��!��/g����������~_�:��/�+@����|4Z-nY�mk���Ceq�}_,aW�e:�m:(`�]�m���#���b�Ee�,K:�\F�S��W��P�z�tbT����DR_���F��]dZM��g�H,@�\�P	'��^6 +��b��i��x����nuT��+�tp�G�u��;xD�#/Z]����M?7	��u����&���0��9�L�]2��C�V�	!�)�b�c{Iaᖷ;����!��D+�N1�iC�ǑN?�)d۬>������uӔ!�tS���y��t�i��A䃰�Xz{~J'?L"}v�-.a �<���5˔��ư5;]4<j5,�5��u����F��Y]��0����#�@bt�Ԣ�[�P*e x���}�Ţ�ځi�k�6��7���C��r�x��5#g��Yp!����Aje@$��7��ATPA)]�z��{���3�X�sgur�E8���h�Hm45N���K�܋�_ެTz�A�%�p�R`?B��X?phq(l�==�OA�m���٥��ݎfxn��(+�3�W�l,�. ��V{>���}a+u^�]��t'�^�}5�fH��sr��|��V��0��̼9������K��7]b�'!o�N�o�Vvܧ���y��M��k p�Z�uE�gIbbrΧ7fy��|�}�)6�Y�?����!L.A�9��k���/�Uc�た�,Ƃ���wk�0£eZ�5&�`.� %g2����h��걐0��˾:���Np3	�|���B�H�I��)	b�Յ��/]���@j��`"��>��]�q���%ސ����ٻe�	��w��~��2���z9��f��
���&-�Imyl��-~ �?�J�v��R��<��"j@�C�$n!�!J֏G�g^н�3";����ĩ
�$����|�{󟔐;�A䃳|Wx���V��J�\�n�fK�mW� �q�%�)	LbEլ"�_���-�{*0�~�x�'��w�\I����
�U�$����e2�5��xk!�Ɣ�Hsh:e(p�!�Q��-�̿*�e�v/%��/)�ƂRw� �IЌ"��R�e��>�]�����(�X�
?8g"�0�gQ+]���� �tFQ��[��20�|�!�`9=�_�i Aa�p>���5�7�����u��>�|9g��Iezg�O�A�:ig5��F�)�وQ`�$���Y*���I�^˧X�i	�×��8m�����
o�ͿDF;{0׃Kz]����/�.��0�.d�����&UHɧrŸ�N�{Mf��4���4��9W�@8B��ЙP��0������%*vA�<+��7п�kZ���\��/n��HS_/
�����+�\�bC��d��K��Ď��@���{�hw�e1��`O��58��|A'�q9�F�6�5:%i�G�$D)�ՀR���L�p69�sI����A7lx!)E�W�:�qa��^'��j/)���������4�����j ^�RP��-~�ЧSNu|?'&۪��S�T����E�M�HK�"�b�D����-~�;kX �Cww�q���HޡNrB����|�W����l�ᔛ���c�^���p�ؿQ�����6T#=��K(�8��������O���(EC>�=�Jj�	(n��� =�%?�,t��˾�F���������o�Z�J*4�9�9���T�L�nBPݢ�Ɔ������p8�@��\��<��ǷO��0��H�<7c7��T>�y~���ͮSO�m���M�zdA�U���:I��ｻ68W�;�����k���>��S��j�0��e:Gw[~��a;?�R-$4c�@�/�r��k|��}u�oN�O��}�<Z����~�j��oR��U"�����$�k�z�Qk�MX�^`9w��:.GMN�ۥG԰~�h�����=6��s=_S��b���%H����p �tꐲ�("�~d�ȄN���>$o��p�E�c�~�!�a��h��M��_i���)B@�����g���.��]��(�3��@�*\H��
a��Ow�G6��궒���^o�)?n5��%Ð�8�d0��]�c%Q��ǆ���ʹ=��Mi����`����0�ld��a��u ?|��v���@o�d��s��j@��m�N�>����J$Y��$��Z�ܖ���;wHr�<8Q��5�ǚ撖�g�^q��j[��mؔ@{·�	G�X7����l��J�����"�eB��@�l�`��V_�7])e�����80m���y��LK�j�4�N�k1U����E�1C%Y{d<�c�Ƒ�����:_�����ȍ� ��G�[��B�/�ܠǡ^��v���4����W�bU���;�)Y7�H��7�7U[;p�~0l�T��&ˣK��W0���ʮ?=��HD�+�͏^rI߄�V�͇��K:�����媨��Y�G���5��,�{��V�E��(Y/>�ho���j���Jjd^��`4��IxM(|��d4�;Qޥ��P�����)����F,��sl	��k��@�o��g�A��e�H�`W
���F�Z3	�o���j,+c�G2]EG������EAz�Tc}>Ž�g��H(�TB:��o�W�U,��j
�lv�sm�>�ۊN��MF���,R<X��]�Ki�}Y��~��!��I{U%�/E6��h�e��o�ʫ-�HS�5"o��\ڃ��abK��P�	HBL1�2�s�;��ئx߄���o���Ӆ�����L�%��O�$kt�D	��'��|&�f9ƜD2*��+>wnYC8l!�_X��l6|J�+��#��K����Z��$>��qY9��O��g��P�ym� �(�F��W-?�nsBe��;f�buo��j1���cQA�mh���̚�����9��/P"p�4�)G����K8�4��"w��oiv_�Ȥ�@ o���R����2��%�`����w���ϰ���:z2x_�ӿ�]B����~�Q�.`�V��S"^T0?]��]�0�䩙WPjr]���h�p���\�D]��l���q�3+jl��ȭk,�ˈ:�,��� ��d��5�7n?:N)��V` ��3W%��{26�R�&i��~y��1j
�J����s�������z��qn�Q�2�嶲�p���>d�`[�+���j��C�5l7���G�\T���׀�"�ջ���m�hr��m�i?�Q]�/����Nz�,Aք�FJ��هr�Wt�������R�4�:� W|�'�d�hCڽ{1F�U�6[?@���ܐ����̓��Vp��4L�==�K��7M$h�����&���뀌��qeJ�����9��i��
�^(�e��zntq�����q�U.�R�L���t|��}^ܭ����z��n��(� W�9�o1+ű��l��L*)�^��c0X��m��Q�@*k V���"�(�=�e,����p��Ƨ��W� ��u�P���o$�����cBh��8�0V]�?�3��|��[�W��G���.w�҉t-k��=�9�-婴����=b�q��t�]P�V�h�sNE�:#��&�y���,�F}�J��p��s�]%@ �=[y��9�>��+b��p`e&�ŝ�ݪ@�yP>��2��A#@�h���U1)��_Ъ��@��*�_�4�������-n#;��/!��6n�-Ln�t�y�:����c=R�PPf��:��.4��{��>r�k&~�~�T�|����`�翔"��TCGQ���������S9E/����o^�еb�vO� ME������2#����?G��s���m}��ݲ㗆-� �`Ea�,�Bnd������C�쮳)k�Bxp��$�G�\@Z�;��L9W1;�eTq ���"�����)�(�}:u>]�3w"� ���A썕�OV6�O\�/)b��P �ĝ�P!f]��Kc�/n�	�,����LkH��=@-W(G`�rl�{�ד}�Fr�^��)�qy%���&��9!q�5��G� ŕ&A!u�\4#����KȦ�g�4�<FE�m,��s˧���oJ������`�ť
�fc�Ca����цZI@����:�r��-�V���Ԩ�b~(��5��+���Ҍ���>r����~�{����s���ks�W��`\�����\���t�=��l.&���k#E�j?�zY��h5�|g�5}�\`Z%R:�[i��uP;���ܜx���[{tn��	���a�]bC�SC��UT��i�V��/��n���eɶ����,�s�V�#�G.`Y�`�zG5�ک�z�ٶM�.�|�õ�C�uC:0�޻'A�fl��˞ԅ$���l�OUd��*g��}�'�pI�مJ�!�h�~�c$��rd.����I����P�q���(H��P(Y�����S^�?]�+�W�V
BEހT�3�Ǭ���N��{$�e�=o��y�D�����y�n��۪����;�9oa�UX����`s�`m>_O�E��T��
.�@0�R�PmB�B^�:u��zG������v�H��n����+�P4�bgd�x�Sӳ	�E��T$<�"�٘���q1��|���j�2��8��C����C��
��8�~�H����R��M��/#����m�Χ���B?k7
Y�W�/kH��!u��S����}�Ռ�AHi�G~�O���S�.��َb������i�$/8?�8������Y7�^�j�8ĝ�z&���ǽޞ<u4��yqy�csl�a3�������֞2\獔�����,�*�����ڑ6J�Ȋ��2O���@n.�HtI�δP�# /	��<sP��ӪV�f�fW������ە�g�b7D1d��;�H�;�o�%5�U�uӤۣ:��5Rt]4���*n��Jp��"�x������V�P=��P��e'5��p��{�<��4�$PlF �B�1�譇z3�&��p/�����L���nspN߮�nK	lYCI�W�<չ9��m$QO��f��a<-�qVtب����h�8N��3���_ي�ӫ*&n��<8{
X`� ��N6����W���#(��-&y�m��J�w��a�BQ ���+�/�i��
���c˒O���d_�|u-�B�������~&���t��#�k_z��`��- ų���.�S,�2s9w$�)��u;�QP9Ⱦ���F��P�9�Q��b�����(�}�/��#7���"2m��n��^�i���Ol �M!ev�%+
jV��E�4I����m@>�N�����*�19n�y&qX0����B�����}@)^K�c���H�\��SL�CV�}�knwG�O�
=<Eg � �S��-r�Sq�B�Ә;ǬIt?L�B����*��c�p>;��D�b�^ �f3�[�K�:0�ƀ�O(T��T^������w+@=��u6�����,� ���m~OgV�죛7K�j�f.���n��	ϝ��%
��H85�.Ķ�|b�
��鋟�Drv-@�S�CBE<~=�A���џ]�|r��u�aPʑ�)���o���?ij{�LET���T���oG��}��.�d.iX/��*�ղ�P�H���nB��~�o�Ү�����,`F�)���<����ȼ�û������=Ń�T/���ﳅ�Z�G8O�������{X-#]�N�6My� ��.H��I� �Ϳ��9����D֯���|�i��0���3{ ����N2���uI�T$p��W�2`)�'��7�1��j(��Ƞ����؄�B�"7��í���|���HϿ2�?2�����W�#���k�a��n�u��ҡ	�Q(��bC�����j$1�!��u�CMp����6�0�8��p�gd�y9e{zj"�ՃCB��J:��n�:�n����.���D�q��KV�����6Q� �����WAռ�	�����m����C�n�`�ҴG�;�?���H�j)U�����\�<�Ͳ�g�4��oIW��G�9I����5#wR-���p'�*t\l�U&��g}*����{"B%r�Ų4A���
�- 3&�d!)7��!�W��*��li�B��r��tl��a��Mƅ�Ȣ�𚔥L@_�V����֊���}!����wix�my�%�)�-c~\}v#�-Xe��5� :���o)�Ɣ֒��Ga%e�G�A?���g�J�uB|�e��ycuJj )ߊ��*,�~���tJՈ�FD¨�!��.�Oa�
�,�$�GMY�Ѓ��u$�Pc]D�K�nEgBV&�����ln�O�sC-U0)+��]�˶N�=�Zh2P���`��?��*�����^!3/����F?�㖌:�Vk?�6�Z]>L���'i�t|�`B~����xs�~M�1=ϱ��/���� F�n�ۍیwh�����~+P���|�t\~H�rvg�bꎸ�P�T*�#�\� ضy,�L�3�h`(A��ι����g}���S���s�qk:b5���!<o�va��Yd'ѕ�)~%�p�|�@<7BD�����~��P�X?��(p�`?-V�9Jf�?K~���:u�,Q
&�q�}�ת�C�)�pŴĖތ��b8�,%��}>��g���nDQ��3}�G
�5��h3H�v��`jf��P����`�n|�])}��b�S����[��� ��D�Ӟ�Wqs�
�*�2?�:Z���nwˀc@�YB��:hR&o!Q�z��ش*��B>�����A�s{�K���B�����]�f�I���k�� �y���k�k����	pI�ng�oy�����r�_ca��l!��L����W�a6'C�V�� �~��˥3(,��Z�9��2��l�@��F�o�!l�[Z(S���"zW�D>�} \���Y;�%i܋�������#T�e?=�K��ia��s?$/%�׬s�?ٵ ����&z�����T.!]�AO8�����V���K�D/�^kK$��v�I$g�Np�������kb�ŇЇ���8v�5���p��f�(W����j�9
#[6,g�^56�x-ֵ�Lm ϸo��R}�> ��mܖ�tm-�o���ă ���S2�J���������9��YVx%��9#�)��Q�OAGo���2G��%s�lڹe=�#b�	�"��n��\�)ބӲ/���FGS�[]�� I>F:�?,>&�t��9w����I̎� Ԁ1\��!|�-�97�B��|�Y!_�\�Bs�4XI�-�;�� @$7���G���ﲺEI��kv(&[�wI�Z+�{��`�ۨk�-<���-3�Ř��/)�CV�`�ci����uQ(ڞ����ᰴn~�h0���B_�Tf����Z8�i��_ު̱ϋ����_o"�y��̴��G�>�pyP��c�k�	$�8؛�(���]����h�l�S��]��e��OX���K��-���� 7r�6�?;�����@�K<hܞ��x	0'�������5�������%G�"�>+y��n(J�.v�ʷ�d��]��<��f��SÀF߲��dx���-E��<����L��	�����z���( �y���s��"cYj��a�6:̑���9����F�_���eN��� �'�m�)�N"�@*DX�9�	'�k[H��k��%�e\�C_6��\Jũ�^��_V�_�E�	�C	��?�ݹ݈ա��H]m���y=d�n��<=l��o�d��ط�u����M_��TY�	j�鐀f��zcyQz�|L�hI� �P"&��\��l1���J_.Y�[M���k%�)�!�"��<1���B��{��48K�fң�J2�}�b׶0h�~��3h���$�쟭�N�8>[S�7��	�������Y�i��%?�u�X�0�
|���Y�N������
�釪�-1IH��AS�C����"i*��� R�C�!���4���</�@��b��r��}XI�=�v}��a�l����A�h?�ZN7=�k�A/(��rZ��,|��S
Z$+����)G�LcOh]F��r�R΄@�M�і����îP�#�4sݩPX�q��og� `���"3�K��t�u$�U-`"�#P�5b����oq|=��i��������>�(�A<�|���� }��s��������A����/�|=��%�;wh���{��ה��G>
o����^�X;ijf�n꒝]VFP��B:�6p+�M]缜ds�7`ǩ�ߺK�l»E1�a ����j�Qo�ԍY�"�ѽ���b�ǳ1#�ۂ�D+��o�Xf�`�v�+��r-���۩�o��}c����j#����&6"�Y��F:�A0��Q��;�'P��e���5Pgq���o��,����mw� �Ꙛ^���-�|��z}���G�D��%&��#��3�u�[����t5�q3^S�z�eB%��璉�)2�Z���3�ta�'qM�r$�ɮ��26�rK4���z�����z�[1�A��y�N���פ��EB��M�zAtyK�E7�P�f� ���-@��g"���/	�?�y�xI����I�� ��eƙ�h��n�ӿ҈��[`x��|Zv���H��B�}�rۆ�����ZsS�N�^�q��p��m7�v�KY����"8�|����*��[�<��U��}�u-�����np�I��i|bd�[�� �vPy�ӹ��-��-�ul�D׸�uMo��� 	��n{�]��=���~n�$ k�AfD�4}��I6�	B;5��������7��=�)�l��04�R{/&$����)#��K�g�$#�M��N�"�CF~�\�cHm�=m�߀�oP���]��w���V��0N� ��ix%���'������6�@�S�K2��'u�	TM��#�ᬐQ=���E�/�,��Kl�8��HJ����B���0<��\�~���{7�cI�����gN K���ϛ.�����4a7x6��ʖң�bK�G��=g��I �:O�ʶ�j �mV��b8�$|��ʴ>�.��1���*Y&��r\����`�ë�~Nqr���	�\���]�7� �_m�o2�]��b�G^/O��D�N��v�ֱ��!褮ժ�%`>��M�8�C��"�����Z"C���+b1,L�;�U!ܝ��cEx�������iߩ�(�����m�N�� xU]�d���Wo֣7r�oN ��,8��O�,ͽe���x�
L×��+���u��+1t�%P�k`=inT���oh64dj:d�X)�:?��8@4�v0�1q�C���EݺU��B3/Zp�GDM�F��	�T�pS]��z���"�l��������?[	XyNJ�k)�w�Pj���g,>�H.im{���Ik?�!E���`���ĠdH[`�?ۧl��m���_D �6�EOt6N"I�o��-G3nF�"�]�8��m/u4 ��}��#e�7 �9�ֶG��m��#\���� kI�Fgj+�n��;(}i�͇��k�l�]�[�����W�K�ċ��!�YPA&��P�'aB�)?�f
f��9Cx��l� ��n�5�����-&܄�|��N� �)E��rd� �%����zF}N�~�&�hM�<�~'Ǆ��0a�#��qb�$w���'��Js�tyb��n��b��`DS��d���M놘n�K/��<�X�%R�9��|�_!�����$�ݹ�����)�ǌ1���{ګ.%	`o�W��P�
9+O0�~/�ZG�b
�r��13<i���_�G�cL�A�,��z8�C��%�����i�r�R�!���H�b�M�k�C^G#Z�fx�Пm�/Sp��|
�J����������U�E��H&J�/�YVp(�(&q�&�����B\��?�-!������;�?���s���gf��+��&��޲��.�W�gz���K�1�}j���ʳ�|~�i��T4i<� �����L�h}�6
��N�m�@��r����r�V1���{(O��L;T�B�]rM�#QQ�`^	:�(�ʄ�o���#�b5%[-R��.����mJq�AX�j�\�Tp�m~�1q���V|}�4�wK�x�u�D�~��h16��G��P$���Q��8��i�qn� dU�[.���#�|����6� ��+��4DF��,����a�m׻1к�D9=�2FþL�������2��HYI����4Xo����Rnx�k����Rk��D�y6�WÅ·�)����;W�v0�h��^>!|7*��7et]�O����?ͬ���h���]�Eh{D	���y��>��˗��D/_*C�:�ا+Sӝ3V������M��f���|��o�k߅a��χsA%��`1���p;o�˓8����Q����-й&D�3�#=b��~��'LO���	
Tt]\����Q��
V�����Nup�4u�}S�#{rd���ۊ%ڧ��[[�?$O��T�G��߽�s��6`����a�%	�%"�@ƭ��V�oaW�m����\�͐ǳ#A!6�0lDL��dk��ubd��*�c)[?�%gURʥP��2C�?m�
���ۆ@L�k�-h�N�i�������E �6�-��C�E�罹)c�R��j�n* O;�o����f(m��Ч^Oϑ�PU��k�픦]�Zd��]G8��<��u�+I'ѭ��uB�N� �FZ����3���#l�o�"�Z��<YN�r
O^��HJjVX�$��J��O;ӡ� 4�����A�Ʊ���9�HH3�_��� F��hD�^�!�5�ލnI�*�sYZ/�v>D��iV	�=C��$5�_D}��3�n��y���].���a�b��������JAl�UQ�O�@��&aM�e�F]�W|pĴ)a[���C^��#oΊ~�|��wa>?���1"��!�w����．����F���ϑ��	ac���h�w� ���B< �܇-�zZهn �}v��\`Z���
��7+��ڍ4S���\7����c�Q�T�D(����g��M�����RH�_U��~V+�{������<V��������2���"�E�@�ǜ�c�KVBr8e�\���(ʨz-��$<���cZ���2�z�G�X�lΖ�����_�����4�1|�2�?���(����~�n�l2�������)ϸ����A���ˆR�£��K�YU��a�2|���%����j5E�������ڟ&��bu/J �(��2� ۭ��o�����s��Q%�W�+Ӵ�yS}ͻ��	=s�Ogj���X�:���� s��:�s����Z�Ep>h;|�����������Ok��&ɠR3]���I[��T�����S9����N�Ӆ���P
��w�y �g�]��Ÿz�k{���սV��lغ�����[��|AZ�F�z��JW���J�~�<9ߛݹ|hm��`yL��`ЯN��I�s�^���ܠ{��+��.�T��O�O�鍨�ʧ0�n5��t��A�ym!�u-������)���Y���$�-��'U�ĺ�}���bA�8A^� �vԁy�W�q�UK��x�����8?������7�K\Y.�Pz�������,R�����%1���
4�v"�[�.��	w�#?�KT)��ʥȎ�i��R��VT��3d|-Ո �����K��Q�����&�`����+1�o�#�!O�]��<��(d\��h���M��B��$琙׎�6j_h�����"R�r�_����]��v4��kǒ�n����-���h��� ˞�*,�󇆎,�z�<�_�c��l�_YO�בz�C�Fɝ��3�r��

�����XAiwވ����[n%����R��q�ǝ��C�_D�c�Kx���5;jآ��wm#�� d�F��E5�R+�_�/9m����T�bT20�tpN����vֲ��Ҧ���?�k>��5Dh�Rג��W��G��!�K(�(��ݙ0,EuV]Z���G���MO��=��A��U#Pp�p":�,f�i�Ҍ���ݼ�"�B��7!�h� ��JMU�s:�F�g����H14�5�xv�R%;.	�q��J�g;)�Q�8�������8[��Vg
��i/\?u�֪~8̙�㻵r��IPZN�*'��0s	?��\�g���Sd��ڕ�^�m�|-DI/yT������n	���� [�6j'��g�b����5���eh�-�'��_�<�ҡ��،��8�x�!O��[W�#,�_�ף5%hT$5/3l��,�����w�@G����H�U۝���p�o� TX�2����E2e[M?p�#��8�۽�Z��Q�R�W��0�_�D�x�$�3"������56|�ZH�03�Q}\�ԌDE)�گ{��Ɠ�W��l�ͱ-��j�a~0}�3R�}�ug�,3�b��`h��Lu�и�6�yy���\�8��i6Ih��7P����M�4ً����16� �?C����(G�ҟ�� <e�Ȣ$��,E��h�U��R ��*������⬚�ƿ��{��.+%D�N�l�#��=Ѹ��y�����1Κ�H�ߓm��ǚ�F����
w3���L"�j�9]>�m�Y} z�\�ɲ\��*��uh���z��V��ԖC��+_:�[��#�/���6�P9�W{���';��g��K9K��;z4EW!�����lmY)鐜��c6;W�ɳ����]�>�}�QKH�,��g�6�e��NѼ&(Z�9Io�Y�JK��8=�1JU�b�<�HQ��y�_C�-���^��S]��C�C�^�V�!\J6R�A��d��D������S'�+�����x�,O�e-�2����(D]4c��_�N�
�)��.�Æ���׆G��Ucw�A�*�����I�7�ƻ�\�(:�o��W��0d&��b��\�O���� u����Z6� ��j\��&_wf+��xIﺆ��9�5]{��V%T�H�<������y�zh2�?�^�e²��<�ص���h����OTF1�
� 9r�KO�fd���0����<+��O��)�k��ʘ2�S���Y��ˡ�`6�pj�A��	)Qg�wi
�"�.�w|�*����U��5�4U�����߽��?��as@6՜�⪱!������q|x�d^�^�	��9����-��9T�����R�v�����4o�������Dy��h�:wHėZ�s2RņKJ��S*����2-�N��������}�|.#P��M2��wǟ�����~�q!���V^��UƋv��ag���T�  �X<)��0!�E���	�|tn�k ��}4ϣ�6�Lx-�u)�����r��SK��B�/3-���M��Qב%��	�����̛|A�"��7s&��$�@슎�ԫs:>�C�����9N(�O�Gb��6�����>��LL��%Cq������)Ӓ��?��?tꌤJ�<!�,��|tLA�nNSO(|)Uaq��n��:r*;c�Ѩg�!Ơ*#.�F�a�����T�(���+�n#����s<��1�ʿ���Z�=�k�z4DBm;�#��W�ձ{�����r��\�nkt{~'�߬az�D��3����͍�"/8�E��q,�A�c<Nqz�P_��1ĉ�^����v�9��\¯k��O��>�M����r�����,w��>�:�3~6��,k����8�����tE���"�2MW�C��Ab��{�(L�}�p�
����+���>V�szX��[��������V�!���x����n�L-1�u��s ��X��['ٹ���X���g��@X���q���Ⱥ�Y`�����P-�����HPFe�,@��`�9�Mc�~U����T�հiY��'�� +�m�۰�4�y�sm�K����1l�7ۦ�=�������9��ks�u�!&���p,�?;/����۱pJkG�W�ļ֭�#�Y:��u=8�w�k�_����(v��PWXR
ƛ�\-�ђA�/����,���EO���}��꽊��%:�Z�A�%m���1b���j��,nsppN�p�wܔ8�^�V,���{)�e�أ|p~`���:�5z�7��gIը��fx/C4yW�"�I����c���f��? ����/<J��1�������w�}��t�ZW��s�.�x��㻣B���ꀮ�o��%Ҋ����Ya��	��V:�|CW��|k���$;�7�(� ]���;�b���i���M��A\�տ1[(���(�(Y|�4^�w|�a�bg0�@C;��|>�}<�B`_e���GF�)<���U����#t��M�������E<��L4i���M7ې���I��f�����{�[��
>�Q�y�����o��bx�Ҝ���K�#�:��M��ù�J����z��-��E<��
�m|���3M������؍�hוb�i�ƾ�`.��h���Z�A� ��K��Sgɵt�>��ͻw����z��-LQ�F. �d���!��L���h�U�P�@Qe¼)9���(Gd|S±��zn�+J��e��`���r�dy"Q�Z�ӅBЏ�w��9��fL��)�	��j*-�����Tb�Z���/�# s��[��,�i�.�3� '�J�_ě�&���^�����L�h�?��_(R�����˄�+n�5Z�e/���Ý��X�n��4SWV��[.|����z�����	K
����d.��z^;�H�3�Q!���T��煝'���rK!�\�s�X1x�� �9tף���v�0� 7�(�9����U�����f��n��8��=���W�F����V����p�.ǰ���W�'ω�I��5?���?���6�v �#|���2FN6$8/�MiC�*�O:bo�Ts��{�������q�7o��>q=ܳ���f
���B����h��F/0+�J4 ��-���|XЫn][��W�����Z]f%a�g���E*1�.D�7�Z�f�DN���?�w�*�P���[�!�+kv?��������y�ӆ湕��Y������D�c����5h�uLl���Rb���u�)�W��n��Z8(�O��k9�_��g$�R�{D@���{�$5��ʂ��@S�涪��9�]��	+k�^{�����è����z&����,�A8��Sppwv�������|D�xCN����dØdG�q�~/+�A�u�º_l�3Ìv�X��
GW�{��nm�1h�m�r~'��"}�	�g�겵z:0<ƼFig����;�m�Pk��AF�5�Y=$K�D���x��E�+{�[|�Ӗ����Z�P�F����ɉ�8�h��7�b�7	��u�$Ox�}��Y�͖����8Ǿ�U8}�@��i]:����Lu��Y��N!���\���-I�pnA�\�_r3'Oٯ��M(w��d�*c�C�z�&�;�o�{��T
7�MB0=�,k�J�z�ύ��c�Q��BE����yfM�4/Y{
��2IF���;�n��G�a�R�]�3�k+�Bk�̉�������s����R�(F�o��Z�^ �
x]���⯢�#۔7��йC.U��/��m9x��9B��T#�lIڹ��sW����ĲW��ܷ�z�=��'�)��?�(F��&��$��� ��X*i%l�,����V�rT[��V�99{e�l��j�׊5���̒�C�a#B$�����%."��w�sa�����E#�s$�hE�AH/�qemK��h��[�G�� X<Ǽ��I�PQTZ�E�~
��&PtX,`&fy�oc����vœ�6�b�KIǳ�<��J������?4
ƥy&�M����KaƼ�(�2d�|?�etXJZ���� �#����F���V�ƿ!`��>B �5�iZE�0B�\�7�-���yT�Ϝ��]/����{Ҟ�CB�04��?��t gS�#f��"|cN:KPi�|N*ЃPl��O���ƃ�sh�ܗ4�|vb#���V�o�$=�z�l*Mh�V �</��'�ـ����٧Lc൩�Y�d������amgc��K'��*NF�x���O��'���({�?��O�ͦ��P�y�~�!��6���`���I	l�@�՗��m����b[�\��,�xF��'��C*Q�՛�oT������hm��i
�>��c�gm��T���� �$�13(i�c�r���|�6k�`�6��_s#������o+�[*�Z�U���}o�A���f�s�e�7��5���n�B��Q�қ��,�7�f'���T�K5vHY�i�����8["դG&�#F�E@��" ��~�UnJ����i'��p��9�^.8��di�����Y~.>--�g}��1J3�u�ܡ'���/&�����v�T���7�_O�X�����L��G.q�
�b���?�6��n�5���r�k��@�%��G5��z	�O�>6E�p�O_2��p��@&f$1��ԃ�6hd�R:�9���]e����ֳ"���/�7#�{Ps����8���9�H$6 Jqك����\�Z��P0q����[6���C�PF
i��@8�Z�\.�Gf�k X��R�&@��`.S{@+4��^��^h-Lwɭ��J,m��0Zp��?���R�4�6��L������j#+�* @�����xNv����J������̴����n_���^�
�J��9l�Etx��v��{�U� h�$2aI<X UqY���y���|��#�<$�S���F�F�����Ѵ34�g
m�D�����.��f7��ᑠS	���@��)��Ҡ
;u8�d*���ϖǐ��I�o�k�f���5�`0:���X���AlG��S���ih�G��ت�W|�I���#�0V/H��$|��s}U�h%;�Gh�F�)`�-���f�M��2�߆%7�`F�΁O�d��kh��h���Ǧ'���,�=���)�5�.�&��?��f_[K�=��"4��'|+�O��12tҊ>߯�ڜ�kZ��M.w�=+q(���h(��f{�u~תƼ,T��X逊��{�� 	Ԑ��zBv�C�U8,�q�&�g���}z"I����$e3�{�
w��"M�|����W�:�־6�?�{9�r�Z���Џ )���<&г����a����3��#el�n��~�G�żJ�ٝc��P#�+~<\ �W�$h�p��D��Ie��J6	%��Ҽc�2�)�o��)	W_��q2�u���N;~1d4�`��4�ls���7�mJ3� �F�W'dr
��a-g[:�����ҜC��B^92�g���!Τ�>�������J�9�E�Bz�rk�pA�#=�(��1��pY��?k�L@@�������+�,����2k���J �
TpQ��@�����փ>������G �~6�?��9 �lO�Tc�~��<� F���J�:�=#�<#��>b|���_!��NK6F�ol��Iq�4Ҩ 3ݝѧ��$)�"w�fkc�o�S7Bo�������꣸+����� J�.P�D=[��mR�"sB�ϋ }����5��F{-ymH�����OX�8 �{�e�t�=TZRZ�Hf<�� �Cb�.�UWIN#�����KC��
Qj�r��ύ/Xg�*�̺�?�=Ֆ�|��w��0�& T>)J,��R��W=��J�/6w����x?5�A^���h6vX�R�<6�|	�#�_����;��r&SKp������ 
9�\��?s3��}[��&6�9�^!QYU�����xFm�KV$�G� �v�|���ݕz���%�/�^�#�w���f�s���v�$��}�󉌺;˛�xQ��*Jwq6����N2�E�p��F�ӻ�I�v�[&n#�%��;H�d�n�3�0����8�#��{�`�J��(�wCrT
�	G�1;����Z��s�]��`h�Y+����6�&E��B���/�U�OW��ۮ$�(�REkp�ԯ���'4f��T`H�b�	�L��u�#p����kɰ�)��P9�+�k��B���<n��l��Su���柿�Pα��.�,��I �����i��1FB�DI��]���?1����|�- �!/G�M�
ß-���R��&�	�%ya��&��a�J`�$�v"�ö1<�;R�S��K��'#N�������0���6>	�H�	��̯s���H�p�mb&MR��}��Y����r�?�h��c�vI��;�� �<�<3�h�ֈ���J���}]@����h�N���Ag7���$���q���U���-X  @���P�5������"ql,·��������1/��dQE���aEذ���</����9}�P�D9^t���G̀��jͷ�^�Z�}@��Y?:�,2��Z��3x����~B5e_��Ge��z�<c��
��l��f�� �v^gR:���3ՙ�U{��LMC�|�{b�R:i0��J�C��JE�@��<�Dߥ��GNr���B25�E������φ�á�R���Qa����J\�M)��Z�U�;��݇+{�$���cNd<jz	�$o����w����	S���؏cڠZ7f�?� �:IlI�M!G�%�߈{�+�����W��y�O0�hX)JyiGw:�@$$�~e������n�*�`�u�á3#��	~�e,4o���� ����S;ttx�0�����{�§g��g�]#WK��g�b��1G����kGA/I��ĵ��[j�gb_�3�+���Ƚ�[8��#]|��5�uNv�u����d)q���Oo�}��JT��nk?$	ꗱz� 4����?濛��5��~BQR��M�I�Q�T��֏��ێ�S7�}�����h���Dw<4�B����V4�ې^
�
��3b ʁ��0��N�-l�ז���ɥ�ɱ)Uvbv�ei�|��\4�z��uJ�D�z��}�o��������̺�QC�E�p�µE�uMj4�BC ~��6�y�?Q[���Y_;%C�A�M4Ja}�@a��T@-�{���W)���8<�1���,9�*�y����ď(@�ݳ���}|Y�ni�$���[����YY*z����^����fI&����p�-���=*�3b9�	���z�%��|�� �{�-�U^�-�	��oɲ�&�@�Z�4���H�B��83bG,Wzy<���96�V�O��s��������#%ۣw�B�L�X�� ��Y��Q�j�u��Y=�s�R��)�rJ�WU=�W���?Ua=��I�a0���\��mg��r8I��u�$�q>
�lF�1[��|��?�}Q�b�^A���P���SfŮ
X�����D�[ J�xO\�b6�r<�$+�1�^�ݍ8vͿ&��RP��+v9�9B�Q%A2 ���y[�IehA#�c�� C��+���M�t;�U�4�y�8s(3Q˵��g�TrT��-�a�Q���t�9�2G��$ݮ�[bG*zXZ�D���eO͞�kݰX">0a�i�vD�&�KQ�l,B��w��~V�aT�l ,ڢ+����
 �1��{g�����G��ZB�9 兙�M��V��Bk&���vڡ���e-���z�ڃ���M����!��IS  �=��ԕ@�MMv�f�hrM�?5.��o�����od^��3� ^PL�.4�ܼ4�&����;GKD1���7깒�qՖ�M��4n}��y����[�鈢�x�|O�6,��R����#��<�DZ���ڴ�t����\��kG�E�房 ҏ|9�i�5������Ă��o�̮͠y��o��?x�#Ø�Y�n��Μ%#��1H �/�{/[7�HDM�o��i����%2+h���?�5$�Kw�!1�X&���MT�Ղ���^!�k'��y�5,�4[l��0�<�9��.9��0���)�B���W��N��X�K)㟇���,��s3�-�v&��˺qN'%Tj�|���oZu�[TZr��=�d�eo;Fba�_K,A�o��@Ş�;U'�(�VT�{��c�#j�u	W6atU��8�7��J�-/6�ȷ����e�ђ�#�E��P"�ݗY%���A���x��|d��-`��'�>l�so֔�������g!��FƊ�d�Z2k�8�J��!�YA�ي~GN��<52̚�''__H�Y[D��&Fw[�t ��aW��D&�Cj�!ڒ�Ģ����`G��Z��Y}���#>Lg.�^#i��.������ ���aV(���hG�@	g�Bt�r鸯��\��� ��Q�%4
<'$ny��<���.B�s@L��4|"28����b��_�
��A�C	ʟ6̦�T�JW"��L��įCJz�k6��krJ
�r��;�)������ %1L�U!keI�(���zPڛS&όj��"�D;�N��(	g-��>tw!�����.el��}ӎq��O�׼6a}SD x�w0W*c�5��n�B��:/�y���4pg��`��#��)T~��Q�5j{W�6�l�<e���uj��H��bV�9W�'U�3Jd���wB�P��'���EVRi���c�1����~Y䉿U�T?K�ق��kMo��;�}�������/CKec2�P�s �|(���ٍ� Sn�p��on�(^w�ɰ����YBN�!� J���E8q�/��m\4�A�_"��ⓞ�/��a��,M��<4-^���*�XUJ�n'ua��;̸�)����d\���58�a�Ky�����dK2M�@U�4�؄��X�z���kKڌ��ϭ�n �3�5�.t��g��;X,7?�M_`y�us�G��h��<����H���u�����#g����u�T6�`n��bIO�;���U�v%ΤU�Ф�+����[��F$��]?��SW����3%�8��-�j]2�L�i^��#�t?v܃�w�l��6T��[<�����vFj���\H
�,1�W��w�Ӄ���0�>O(��|�`���+���-4�h�	�]`¡qOB.��!��:����6�z��i�����~]:���QA0�/���X�ץ�)G
�;l*��/�OvjJ}8�@�I��������V0_Bģ���pi�$��Yb�2H�3���pU���<��6C����-(�Ǣ��,"��O�X��	S�z�/�5g���`K�à�&�B�t��~���s:_D��sC�*"�<��j���}�����u�rHV�CFh@�u�T��@�j�o�&A�����3sA��t�%�m
 $v�f �����Y� =C��)Ki�x�'�kِ���'�{o4g�04j>z?Q��L�6�Jf����{��x�'G�Z��<�v+=0k�T�h6������� 3bq�t�3N$��l�l�w�������|*����Ն��j����YY���b�L�:�q�V��oojJ�Օ�l7k��΍l�A�c����6�~4�.PD�S�7|6wm4��3.bZ���y�P���D�&�Y��o���_��)�<:�J)�*3���K�*GC�+1OJ�2)."��w�e�>M��2Q��Ec�ᖡ���vc8u�U�U짾�R���h��0%���wU��p��IZ�>��"�Xs�~Yf(r��lQP~8CF`l���6j���$E��4(��'�L��[���޸%�T�)�(#��=yڰ�30�R���l@�像/����U��
�<�I,���5{*�3�I�&�<���Y��ޟb#	�0"0K�s}`�_�g%�Gƈ�d�Ď.FKӯ>3�b[�ǨNԞ�<��������ʆ,Vw�G����xH�V	BE�J���L�׫-
�WB�y*��a����8��l��a�*�Ml;�}b��=4:�G=6�x1������3r66s�t=��Th f�t�/f<b!��Ѧ/�zrC��ڲ�Bk �*��.������n�]�W~��\D��d��\6��0���W���p]e�:� �ޫ��@��)�~���u,���;�Inb�0�s�� v�/�lw������|f�5��7Z9�cM��Ellm'/�\���Вo3�sğћ�?)%  �Am����:o��&�r�v<�xSW��;[�p����Ĳ�!��
��;|�gblx������0�.R��㸕1�5�;>0����sƷ�؆k�D6�}jye�S�#�
�[�Ǜ׍�ωA��s�[�n[��������۲wc���j�WH�8��u�	e����j�Ho���0�`�dm�P�ֹ��^�/ʏ���)�O�}���˅+���z��O��r���������$ԅ�}͓[�ڪU����D�,�#�ߺ�2�i�uj���S ��?P�]��UC��a.�����2�u�_3k_��Y���9���h�A�Zj��N-ͨ�8R��5��uT��)�G���7������τ��jhΛ�v�l<�H	[��dy�ev]և�����l1�M�n�Y2@ATṘ��P
�����rKeܯ	��tA	�� ���LT� s���P��!F��_��w�b	�q�A��ϊ��w(UO��o�gv��d��(��W��V������Û|*�\�)���6æW����)��I_������3�uv �� �
,è�h ڸ9%�l)��\:=o����HX,3 ?����k~覘J k�	��V{���������?��T����~����g#D]����� V���	5Na*���f�zцދ�!�K�x���#p�q�Qh���v���a	�'h�~�	@��َ�r��$�#L�&�P�ݼ(T8���F�DvU���-9��������$r�l�fԣ��')=�f�ӎ�0�,[D�2��h���*3Q"2/"vQvx��?�/�;�b]r���?�
\s�ﯳ6�A1�v�J���Β�?M��=cʸ�Y��Y��i�\3 ~���huCd_p���	��M��< `8����9~�?5��-�ׅ)v�,V2�A�9��aR��𴠚@{v�g���n��W�6ku����L���T{T�w��d�b�p,-��Z�_yY�6(�ov�H���ȶ ��4
��3ֲ�LŻWU�0�X�u�=���҈Vrf^>-�O%��;�6����e� �:�{{04�g2�?���z���٫�o/��P����^@N��%p���?nEu^(�����[xo{����;P`�ゞ�]��}�����:��:���6���y��k|ރ�K1���8Q�g�C�خ	$� P��C���j;~H2 R��]��~�vW7~���������^ʻ�Mx��1]��[A�@���(�P�/_���0a5�(�(\U��YH��S������۞{��)uEd�N��Q��	�]۝��y�)镖h�����+��m���8�����@��13�U�.�/�{�+��ޜѭr�N)� x��b��kk�v<����$n4	.G�LD]��XJ'i�U�Y�京k?d���u�Ђz.>v�o	b�{��K��_�@Ω��oM�M���V��F�C *֣�>�7�:�9�c4��5P�L'�v�����,���a�_ws�A�qҶT9@��,J�sAb���ࢁ�)�3>��~�����甽�$wZ�g7	E�(F�z�QX�;fl�9��$��'z���qBs����Kl�~G���uT�V��/�����Ʌ��o��l��^W�3ǟ8���Y
P�R��7�I�xn8�w�����=�CF�fg��@/�[~Pt��nسcL�����D���Ȥɶo�;����9/��;n�6(B�(^Lۓu%�jIhUzk+AK¯L��H��d�q%M�g���	�A�*��%,?E�ny��;����w�N$z�U ��ݷ.�Ps�o��iy�(�ӵ������L�;���Q���,��+ʱ�}��N�ls1�=M�������;�%�����9���w�|巗7S�M��@���M�k���^S�m�Ue����I5��g���bP�\�Wj\�f��`�F7F�V.�W��ECrr� �����co����[�p��v�/��1����{��{�7! t��b�.`7�ӄ��?����w7��ܤ轱��	`1b��K��n򈹐�]���E��\^{�W�¿�o�{��ERb�J����MaFZlA�2w8fD~UM����օ��e*�H�4_	��xDg��O��C�:w�C��؀-��}l^�U	����ʖm���+�����i��L�0v�p�3�_�D�����|n���VtR�D���m�I�z��jd�R�*`�����A�5%��ȴ q���z����)��^)���8�RH��J�Eh�jЋ�jy�QK�^�5!>gN�|-㮙�fz3l~z�bѦ��� B9Pu�w*�*#���qҖ#�P\�9�xm(
]���V���4 }��MR��G���6�]�o9���Ld�ľ�xi|+��� �}�� xqgn�ON���#��|����K��6�w����a�2Jy	������;�4���-�IzR��L�m4�80� ~-�G5��|"9s��Yq�+����Ɓ=�d�KK�����A�Џ��N��a�y���/�ʄ��/���g��{+����@�����贳<Аr�T�u���/$Q�v
��� 7f�.���
�Б�P�D��ص�MN0~S���d�y��d��t��,7���%g��1ɴ�F����CJl	AǒC��A�&�d� �k�G�=�wt���{=:�z�)@|��A�3Ģ��9�,��a�E����T(͖�N������ed��c��}]�׍H�j�[����~		��~��i�0]�	��Ez36�-�V!�u��HܕH� Ս�Ԩ
fe?rr�:XTg?�[vn���}(��B�@��x��m �$��Ӫ#-�eL�ܯ��,�'��oD��X0�;��DL�j�N����d�ĩ��,�֍�4����HmD`хO�l����ZI��me���w�s���y��qi^uz8�����5��䈜G�ﱿ��.�>��ZYhV�J���Hru�y����N�kבz���^P���Z�+���2�r^�'|�ľ77|���$���~i������	$�M�ʕQ���▒	Aj���H�?�
i>�~@N�c��(�G�����'�|'e�d�
��Q��9u#��*���[��Z��S�]�kE
��_�%H�n���� 1i�Ϡߝ]�O?4w�qQ6��V���g���h0�qH뱬}1��.���
���	p�*�\(e�$V�éVO�)Ot�E��RR'gq�i�S�꼁,ڠ����D���4|&nQ�N���y�U�u�p�J��O�phoB�/��-���;^������8=�av�kC-�(+��H(�*ĳ�����62	�E��C<qU�O�Ǖ~��H��]�=�\��3��]�T��#{ k)���y�'���}HǑQZ���]���.G�Ү�ѷ�V�\!dٶ�[E���Z�j��=���f����g|�W���3����A}NkLR"�&�@w ��6� �%�J��0����^1B�g����Ǯ~Ã �=��R@�^gb3}`���;Қ�%�:�X5c�p&-g���������E;��ѯêa_��w��ռ�b�c�<��u#5V#�PqF�t݋����F$��*�c&<�&Ns�5@������V�@��(5KVT���Ut�����{G+)�@'����o��LS�dmWnƒ.E���>o0��)��g�����Uu�Rk�tw���K����\\��v8����ogd����������ʜ��S��UEDCת]:2h&�����y#:ȗ���1U�z/}}��9�46�7�@|)f�x�J�شG�x���D]p�E�!H�`��K"f�rk|<�{�1*�@�3t��|S��{c�50V�=�ص_���Z;(=��6� �@�:�9�rU�9�m��@�ʍ��2p�g~E�d��@r��ޜ=�{�P�=��k�_6�Aqk�hU��H����[h y����" c��`j�C�y�PV@�%oZ�7��m�C�;��=6� Ip��S(�ڡW�J�w�{c�2w��G��_�a�-��)P[�W7���'�2�$h�W�����}#̨��%��T6��x�N�w[���Px^cx�/�bsbB�Zh��>P!��~����V'!�_B�Z|	�� �oݜ]���"ɨ�fj��Poݫ%P�P��&eb�ݹI$�R�G�WO
�!*�D'�u�2@ ��}a��B�`��c���-���e����<�8�<�����3�w]Z����Q���3�C�2��U9������\��eN��X�6z�		}���Vj�貯>8���� �ɣl��3�3=����/��X� �y}<<��<�S�D���KZ$��� �ߨz"�����_�����g���Z<�>{E����N�ȆaC$&��Y����a,�Y}����
dc��<u����c�����������c�c,;�Z	U�G�k�i��5Ŵ���Nz;��<�x)���}��,	�/��ʃ6%����x#����G��\F���0���BV������3��)K!�����w��Q���1�$��9Q���b�^�..H8�uk�O%5�ꈵ�I:�B@�G����"����5t��\�#Rٚ{Hẑ�����G��W��N\e<Q� ��9j�Am��) �QR`�EkڍqL)vص�Ҳ"Q��=��ކ-�j�=)x��4ɫƀ*2�XI�KI���(�j��(��b�-��ӆ��҉�)�0�\Wb�Ӆ��`�eҥ�,]����.Yl�t���P��~m-:܄�>wk
ˣ�kT��pE�x.�4߀3(�|�}� ]b�m"�wu��.wl+)���d���N�o�j��e�0S�H�-!Ч5����$h:pa�M�ǐ����*uJ��.	jg}X�s�ǕW�_G�Z�%p8�N����u��,����"_cM)O�Iv4r��tfHz���9�i�YM�57I�E�*|m�ǁ�0]��6��r���3�4\�L)�ć{j����rC�EZz�'��֗�D�n�8�q�d�A�k�����[�A%���s|y��[��p3�dĻ�H��b��A/Zj;m�̥j�f�����Ww,��3Q7�TWA����T��ŵ4�={����`F�6����5n��`{R`>�h�=���$�4��پ�F��c��E���X�lj"�-�`o�d�+
oR��a�?ej(j�O�9�g�}�Aj8�K�=>�Y6t��/z9Ë�F�y6C_�z�~�I�E2��35��\��%|숉��熖�ɮiu�(y��
��	B�,����g�O�+[R�,qK=G�e�vx�L�2�h����E�2�m�˪C��yͦ-
Ɏ7Â��Ȕ�:���'�d~��V�s��t;��y0���@D��Fi�&=�4���b|����^딙����,B~��>	KF½��� �B����c{۵q�J\�ma
g�Ii`��ҝx:��y,�_��#�ҹO��*�g;د����n���J4�?��#GoN��h��Π1��x�O;���]!�·t���c2�4F��o�A���L��BO�%/�Zs�8@ۚ���ejw`M"�����$׍���B:���jݚhnU��3]w&�5U�B/�����[�x��=�E���k:��f����f/�hw%���*m�Q�y��	�?�dP�w���QD-�-���N��}��6��:ͥ���� ���cw1a�MT��._�OsN�R�RZ�2y��c�K��!��ûB<gK�{��t_�L�B�<.��y������0b�L�����F�Ȗ�m�eq�����'������/Csu����/m������9Ty#�]g�=�"L1*$b��3
`@(�ƹ�֥.�c(;��@�<L��r>�ʉ#�	mDG��/����2�ndh��E٧��A��p�ڙ������<�<$wqÔ�l�6 J)���=��oE��[)x�2�5 q�q���W�P�J�P��3E.z�H�]�A���0x?c'YRJ\]h����vT�\�<4���q;�8O۠@���%!�e��8?���z}M0�yx��#OG�>"yh2��ɑ���p}٢K�c� Dճ�����GK�����`�|-�'!�i���~|ř�����Zm��е�w��7{����c(��^��<Y����XO�5�{s�=�c��тM����ND���2,�d���X8�YP��f�Tv�L�d���2Ǿq,n:���@՟�K��}�|q]���MC�u���?(��Q~�Q/��
Hs��~�0���~���&0�<�}�̦m�ɋ��`�(��Y�����*��Ȇ��h��TG�˕�%s�fL�&��s����_Ry��س���&{���a�N�s�_�	����;�D��߲�po er8j��%�d-����L��A��|����K�)��P}����J�G��������"�u���(~'\���e֌�W�R���2�
�I��x������=-hk�S�r�;&I�M_�3	�QLղ╜m�Ƥ$�<[Z�R��K�l$ܷ�o_:�Z�%����fXQ�#-�	��B�˹[��q-8��B-:�>��za��g��3~�u�NKL:�آ
Шvm
����1u�e��RR�-P!IdĔu�H�G��	�l���,,��N� �xC6E@u�й��<C�P��_2�R����%SH���rW���xC&6|�h��� �c�`6B�%�]]7�s@5����.M�n�d�H��0&VVY�WPn�$� /������4�{��p�dq��+!���JV��oW��A�@���u)��^���Ac��Z�u�'�}��iuTv��u����x�Zn!E�y�"�
�II��,�Cif��9Lu�om��;Kn�\8�n�ڝ�$��P��b="`|��n�|h��/:��ps�7� -A�@�@���E��5#��A�d#|%}�x��|3���@l�~���UZhH^�Rz5(z�^Z�ݰ�~��E���$�9&�*���j�\q�) {*U�7�O�:5�PO�;bʄϰYH�-Q��u�'�`gc#%G�I(���W��a��>J�U��ũg�>���ұ����yn�\�kK�A��� �����թ�tx�}%-)�D���g���dx�(���^jJE��`�9^-��O1��Z�{���5�zV[G�)S����SE�I�I������:
d��s�����{B�T68n�����bF2
Pػ
��VC�&;��:�2��lMn�^-��e@���x�2�	T�b���ؤxL(ڒ-����[�t�HR�l���+����*���.(�����-��Ը����Q�� A|�H�t>�D�
ￇرr�,�Q�� ���1p=%yZ��zj˫��Wy��[����r0FCL����Y=3��������η��}֚����[~�%�(G�f/�T�;C��ĖM��4�|]�0�V`�	9 !�gC�"�to�,TԀ��㫃;�`A)_Ӳ|��'��dW+�ThD"��p9�,��u����]r)(�7N�/A/ '�B?Mvl���}eo�ۚ3���ݛ�����'�!��{I >YL��W(�en	��"̞R~̃(=�2��8^��`��@0<V� +�М�O��|j�i�s�h�t�E�Tj񖀂e�0E�BU&��H�y�%�ww���C~��Ļ�`��nWJ��U=&Tq�Ó����B$+N��Ɋ�C��#�hu	���kH�%�:�ۢ� ��*c�J��Rˆ!�א�{&�r����f��xġ���"H��U'PȍqS�B�dpa�5+~FO����h����Ͳ&k��4K��S�:L��j�І��x�Ɠ_�|��._�ߎH�!�-U%��q��O�oD�jҼr�T�iq�r_!���R��`V`{����y��4�i���#���2���~@���^��Z��Ҁ�i~e�H,m�ZAK�_���S�=@���>7�Ρ<��%@ P�w���R�ڙ$5O���`�Q�'EÍT:�or��f��S�$�r����/��L�}4ӈm��:ddG��Q6�/*�u���
n��������q]��d���-L�Ov=_�� ��9�c���+B���tϸvགྷ'��Qz��G�B��#k2L�d�8���I }�F|��E�^�~����N/Pv��ĴR����8��1b�snb������\W�z>�_�ȭo#Ť��jȤ3�"2�+ �kS��C��Cn�٘�4��l�n��|�Q��Q����ȋ��E^�D$/�#�4Xژ��m��ڴ��9M�XN����1N7�OoY�v �j�z�2��C����f�[��,�l ���6�Tf��/a���L��7b��=@�5ltx����C>/��H��*���ϸg&9�y؎�3�b�M�7��݆1f��o�b`���TYA�诂w���,%B�������V20���MN>��n�}P��f�z!V9���q$��?���m3������h撏�h/�� �z�Q�93e!aP�4�����k�5��� l�˶V���[_������
:-}
�)�lU�ƴp�b�q?�s�i��?��
[�aria�8��v?��"_I����Or�m�|H��b�BnKb�ۂMsX��M�����z�c��E���)5�4[��70� �E�3��	�4����e�+T�v3	��q���K�i�.��)5��0��(h5*ԁ�%��p�������W/��X�6x�_c.ݶ,mV�2���n�FUPj�Ӫ�2hա��M��>���o��UY;�\�W���[�gWn2���}�P��I�6��+,��U�i��8|"oMu�8��+���(x�ZK�;?~�u3F�]'�}�w�8s�<�f*9��eyM@���sF�:O��^��ɴ�0�h��k���8�b��w�q>����?�g�uwu�w��S��% ����κ�8rq�t�ؒlif�F+"iH����3���������f�U4�(� ���/�.\��]���QyW��d����|� z--?��n�?�61)�W��x���&��Ϻ`$BQjӨN��@�ʄ�^OKxVW��'��qs�\j���qF�{�ml����B�_˳�e��{u���������rpCT�8	d�U�Nа�~��Z)�O���}�b��*Q7�dd5>-i�sL���1���S�j�:c�8-��*�x-HS=dEG���df�ū�U>e���W�5�ĵ��R���Q���+���1�sˌ��uH�nWp��Z��{5���Yh4������!�3�q�[Ѹ�t|;DN[JnHt�&��F3��BQax�U�� 6�(O?,���bd��lA;�"uw�㽂:��ձ�KX:?ZvNEl0���P7�c�����g2�b~]�ڣ�0o(
vq�i�&W2@�T��7�ڌQ<�b>EJ��٘˶��s�����������s�ϿI1��^_?��t��[���ʭ�,I�D�G]��ޑ�j�k��Z�ű���0ߏr���j��<�T�X����+��	����)�o����M��'A��9���0`�?e�l�P"��V�a=;���G�{���1|����/qd!�d�� ��T��E��[T5��Df�ܑ%�G����ş�<)蠝�;���װq��u�L��J��E�:!��V����͚(����n>ʼ6qh3�U�a���hR 6#N�C��騋p"�{��Η��W��H��t�_8o�e�;W����E��VI=M��ߜ�ՄN�!�lH:71��g�J���+?�>�v�3ןx�]�b�pW�o�C ��T�#{���3�K!�b.(L�>n�\��2�I�$@e~��+^]H�h���Ă���0W�Ԅ���\U�b{,���WCZ��|'�[����^3�IwJ����1JχA��ĺY�|A1�<'����+���k��j����ɹ;���fQ�tw������2�߆��Q{��J7����WSC����qJW֜��oA ڡ�h��j�����}M�T�c[�&���¨�w��o��B.�^U�a�����=4�+Y�e�ᤔV骳ۆx�j�?����J��!�eM��S�gD�04�Q�sz��ߛ?�,������-��J�9���vp�������	l ��'��u�L��'\����*R�^�Щ�ޥ�3YYc�E�A�����&x!�l|�۠�p0�� �g���Ғ�hOJ]���[=���ɬ��L��#L� ��M�0��W9�"z�?8����h�}��e�M�-�n{�0�z�l���~���Y1����B�iՙ������ޯ޼�k���zW�F���n��}�L��LD����h�f�+޻6-K�&�S%��a��4�:���{��j��{���i�c���l�9A�%�ꚩ:���i7�g��1��p0��KW�oҸ��1�5&��]t_������ݢ�N}7��]Z>���+�Z���R&�B����LIO�
%��&�g��-�� �vj;�b��f ��C�R�J3�sc��T�cw�E�{�h���|E��u�X�����>��8���b]���R{��ؼ���$bS�Pi��`%[0��3����g	��<wSL�J <�\���]},�N��G��S1�>�I����dM+���Ѽ�&�9k����K�u�_�B�խ�S֞lǖ�/FӲ2�8�P@x��X�F��i\Z�澥����fOƯdh�����=#�F��9cwVR��=[BצjB�c����#�/%��I�?Z�3!��[F�b�&�����,K+���2�J/o;$�B�5ϠT�i�J��Q<��70�m�I�I���r��ܖsiQ���ܲ�Y
�5�tq�kՆ�DAVW��i)�.`�������yi��N+q�ށ*e�T���}�n��S��?$aï���iIe��Z�b�|���>
�(��YѸۀ���7i�q�q�-�	6Tl:_�F�O�L������ {h�>0����ηj�ٽstǪS��s��?���
�xz5b$�6I������� ��c��	�L�J<=P�4���}E|:vI�+�k-WQ�4%��۲�~��^�'�j�D[݈U�3�n?)`n�r�G�Ѡ�{숃1G�������a�Y���[��� �0��,�f�{
z�X5f���.ѿ�����mbN�������f�.�d)�N2 >Dg��D4:��D$�9Ƒ�HCmf�CЗ��};����N!���Dw����$u�"2Ȕ������*Z����%[r'Hd�b5�f-�n(
�يp�]��+:����Y��v�}��k��'Pvb.'t���8]�4���s���konh��3~�tђ��g������3H�����F��ǯ4�;)����J~K��e�4"�:o��~��R�J�X�n'ڥ��<��i�]#	iqY���l|JÍ*^7�
�N2��9�T������d������!���IG"��I}�E��~�ϖ3�~��	��+�sB'[%@�#�� 1y9�6E�l�MuT��"�BCDx��#�q�\/|�NL	6�`xRSm]m;���33��
Y��ǭ.�,�A^C^�/�uM�"L�����:��/���-��8;LD�c^�'�|�
��;e�Q��6Vl�&.}���A	I	(�϶�R$�͸߽IP���+���j�8`�)�>G����y�s�[k�;M��-�����	�Y
d��0Æ\9�(��s����_Y��7���Z���b"�m͗����v�#�F�=V4Ik��Y��Ɗ�I����hg�o�/�b
F	\{dN�څ��̋
5�&6r�����ZG�bL�������:��4s��]�_�M2�� ��kf����z�[Z�xڗ+���\V~Č���:�}^�ɾ@iE�+T��A
+��#�����ȅ/�b%$�"P��	S���w�Z��,��DI��Q�D��oM8�@e���8Q���ԛxN�Q��Il�^!�h$e�����"�įd/f�76�NpFjh��]��8h��1�xZ�iP��NsyF/��0�ߤ�^���ş7^��9��ʒP՚ӕ@/U�mcҽqPwٛ���̇�@�;r)�ʒ��14X	 :�
5�n-���)/�������}����z���o��a˾�0�]%6��=�ӫnJ+R���Q��H��T�5����,����c:��.�S�i���GD����,@GKѯ�/�v�,^��m��.���Ma�=��ڰ�o?w)��"�V�M� 0�ĸ�I�dp�i�c`("�:}���M%f�t���^v�R�5��33غY?��U�wUc�$��)e
X�O>��h̖ʚ44O��(�i�?�qi��cR�H�=�(LW��s��}M���8�^q��d�o��Ng����0�U�����Î�K�#�PTC��mf�"i�UyL�IV�F����;^`�@雸L�X��/��L��!g<!�Z�g5�6Dǎ�iػ)P�MX���V{4u�G�2�BP�!�ߏ�,���}ab^7EYK3O"&V�	�j�����'����+����]Սy;�My(<l���|:s����M�~��@ډ�Q��ʌ }i%�IU��I�
 zIb�ٍBD���oO����^�Ć�r�GţJS��>��" �61n�y��z��c3ޑ��i��ؕ,�8P���E��]�hb��4n��y�
�3{ʦp6��.h=�4�2�`���Mw��M6˯r���~�Z��=	������a2@6�+�^�T3�o�Ko���j��\�'}������-H�C��c-BO�Ԇ<UA�xj���R'#�����x�_&���P]���U+A���Ww��$is���H����{���Z��]d�v�+lN�ecX5�#��O�?�0�D�^Jl`��mY�7��'4�8�f͢gƆ~�D� \hH�3�o�������_F$��}J�v�ZʵI �i�-�Ir������0:�*}�f�){�M�Y�p�̙n��E3���x,OgY�Rxt�S�B�Y�G�ļR�N����i�\��U(�&���yH�?~�j��/�EC<�m_S����]S����Õ��n��5����_bo!�G.G,����u���/����3���b=k�.e��Ow]�r��m��w� �`��D�x�/o��f�=���x85(t+|4"���_[u�E�Q��j�VAm
-rT�B2f��1�5�ev2 �aW��R��	L�.2��V8��3�}w�B��-rw6����g 7��3���5/*�S&��X�U� �>��9�=�q��](M�c3����i3L��9�J��c�����^���vM"6t�vN�
	lpET��:D�ɗ�!���6����P�R�h\P��)O���n.(�t�	���4]6��2-�=X���M��+"t��ׁZ�d� #�3�<1� �=�i�ͳ�H���%b�F�K�uL2I�#�#�z�mZ��X:�x��8��
6%��c�b�����^.[�^��� ��aBQ_�IZ��:��M�C)���%@���5y��F��J�R�"gGm;����M�����Z9�G����*�:~ųM����&�ԃ���g.��F�+���[��ʴ{5'+(�JX�Bi�, ���{w2;m�h��O5O�_�h���R�&0�e�:��c5iT��5ֺ�����S���y����}�̦�9qo�[�22.AY�s����Pw�Fퟬ:a�"�{Z�J�С��ǋ>���/�s/%f3�>��3/��D�-W"����H��bן���T.SŶ�~��^��<c�#��zv
�&Y����%�^�9�]2a�9�|p!f��݈�o���9g��-��5{�$͎��n-&� ��W��jp�:�Ry@,j��M��{	�X@��9.Ǥ����Im0���쫱P�_�����ۗ�̈́�`�h��]|�PBtr\ߣ%fKB4/i�4��wE��a�1�;���.����wV��G�Xp8��UX�wW�\O`���e��Aǎ,���R�P��_�4B��Ě՞�8�GȪ �Z�0��O2�Qtя=;�Z�Bn1oo����g1���F)�X�U��>AG�x}�p�Kx�u�'���`����ǳ��L��~֘
���?�6R͟��Ю��-#,���a�-�-�����s�~S�+���Ց��g�? 9��t���n�1 E�����m�o�Aen�z��mc�Cܘ<w
L�jb��s��Q���`�z
�b��'{���aG�I��im�闼���8�����n�eӇ���Qߢ�'��Ɇ��vQ*���t ����͕��8�s\����$�jp�w�ݪ|�d�$�0��k�&��,�� J�f`k¦�q󐟐���-,^=��wu�ײ���$����|3d��'b���tM�7ZL+.����'��/{C���'s.�쟓	NSVC�6:�u�4�ý$e_T�p:��xHO����������aƺk�8U�N�L'�ӌ⩉>��L�e�O��z��{Џ�)�cQT�Cs�u��Q��El���Zt�ݔe���l���QC�j���F���T^�\�?#�2팤��
�A��,��י]�Rk}w�ϲ��S6�}��/o�r\��*��C������H.M�:1��5l.|�r��!�Afg7z��\Km�zĵ��s��K���%��7�]�#J�}�P��DL�䤜���z y������$� 5G�$���̪��N��]9Y�?ë��Z�
�fٯ�=� �~��:�9����YwX�[l�i�����#I>j�2t�m�B�K�#YO�ɴ@�ӫ�cxg��	 ��.seD�ñ*:�����U�u�o!X����*w�CC���V�"�n7� ����b�,_���~)wMtU�9��� �H�����ݪ��e����B*�A��Y��U�F@�KP����"gv����u�� %��$]m�n_�:�}C�%kt������-6v���4Z�O�p(�4[sD�˰�q������F�����cD�]b��WE����ːV%�����?�6�n�I��E���{����o�2����_	g��qH�zO�ݞ���)�n��F%��N��;�o���ı|���z�R�S�f��?�4�<-'�����(n���ڀ��$����꾺�b��]c�j��?�W{���n��طA���A#�2a/�sa��.6�Q	k	��h]���g̼��A處��:�͆�h �YQ���Q��c���vP�&#'A��>y�_Y�}�/Pؠ�9R� ��v�7��b��b �N�p�6���ͩ,�� e��
BU�N���73�����aY^�w-�a�[BI8} ��l�&P'�y����.\�1�9�T0�w�=i���b/G����v.��0>ׇ����Q��+���3EW��4ċ��������I���}7��=�0h"�$k�l���'Ym���eK��K6��"�[�J�g�o E۞������ܓ�*]3Cu��t}���	��g�<6A�!5oR����'���VӞ��rvz���}s��e�FUH��"p�g�/����y5Y=����]Mr�dBٮ'='^Ϟ+I|�ʡ\��]��d������*~cŕ�t���D<!�b��l�]]~�����
��cw�	Wk�A���t�U"+�[�������I~^��yxw�!�SO��|:g�a�Oyu�4�7�7I�x�tt�1܇��o�
^]����X���R���Ąm~-
<\ی�y�.�" ��#���K��x�2EG� ���)�uLH�Apel	��ۢɧaQxml�ͨ�ϛ��d,�p!J_d�h��ij��{�Н�,��8a/b[��(
�E�m[�@
��L�Ҳ����8����.���P?2�Y̄Óz?Uk  ȳ���ǯZ�8���r�$*�&��+VbOM�42\+pJ{X&Rr-N^�6�,��X�#2��Z��>#QO=�q'�X�����Va^�C��cH/gKRl�U�\��Ky*m�c���9���>`�1c�p��y��D9����.VJ���f#�K<��
C��_�^	�Ӈ����gPg�U�Uk�M��/o���۷:�'\,T�Ɩ�� �#&�g���K�RT�:������YH�جے��N=Q�(ho����$:��,':�q�(� 3f&��gJ��$��NW�道���|z��݂��<A��@�c��.��Z�DF���.��<�YB��0h	~*��g�G_ ����~-�}��D�[b���Ω�����Z��z�<��n����l.�v?�2*�f�k��A vl*nV���{�>�o��1B�iK���i~��~?�eq��m}wD�)[�{�7�����c�z8^z`�2aHYۏ��qarT V��'	,��ꯍ����&�8��q�M�u�]�Y�%��eP�4������n��5��fTkÃ̲-�˰�������'��F[�f ��D0ĸ/���ws�
 ��őp�PF��f'`1�9
L���Os�^q����?�G�Hx��Uo��e V^� 9��hz����x�٪?�G���B���`��^�X��ú����!������Z�����2Z�0�<2������9,c,F��ք�㣻O�y����C���p�ƁtԄ��K v�/\�G)���Yur�n`�W+dњ�U�_{��j�0t���)�F�wr���Pឫi������B���/��(�@Z[V���ʅ_Sp���� �r�([�6��jK���w)�8R��]l�а۔���*�R��T�B`<��p�4_%�45�{>���K��4*��]c������o�YOS���{�:x�|i\���Y�Vl5)R�~��^�}�͏������X�S�Ϗ�q�ȍ�'����QKT3RY�DK�0�5�II\�δ��U\nž>�Ȏ$�c���
��P���ͮB��0ڐH�C,.���]���Q�oî��X��v�� " ��� ����2_�0��cK�2�yb��ˀL�Æ�����;�y�m.#RX^{�n���}		r!~�h��e�4d����]�H����#[9O7m�l�1�+�6�H�5��Vg�[FRɭ�U�7ğ�#��y)R9�oKժ7.<wi��Aw݄��IQ0��Y_�����O/-�'w���A�p��_�	2ˍ�5ϩ�G
|��)+_�E������:��XT�U��V�^�����/EB���=6Ȣ,�h��|�,S��v'��2_����]�"��x�\I�e�V.e�b��>f���r�%�e'�(�``C�g[���tY`�Ʋ�
2$�hNT����4�t5Հ��������VȊs����,�]R�;l~�#�2�F���"�b^a����./���5�a�=�3�P"�Jp��(�-����F���0&��7CY �9�ٱݽ��"�]���g�it�0��#�=y�^U��x��ǿo-5Wp�J��Wΐ���\�Y���yf��w���l�w<��5��"��fR�\� ;�!Basv��K���0��{t����uw��6��#(��v����nw�Q�O0�ya�h{�-���£��%��u���8�C�*�7��8Km��}?���mG �s1�!����ׯ;$툽f����!�9���\L�%�H�f�G�x��<tLb�u8����9_v�k�䙦��y%�Q^�<�� �F7���x2���Ս�M��D�ίg*�3q�42s.81R]:b�G�6.���
ܭp�~�N�^� '9������;�p��Us�_z�\fhi��c�J�Xr��e�a1f)���f�Q�ku�1��<`
^�Y���<��4�d����Ҋ. <(	���4��$�/�:�k��e�v��mp���������5<�p�Xo�)���ʪ*jO���q���˴P֖\2s�d㈑�������^�!*�����:x �JcX�����=��B�%�M���m͑u�d�˭�j<yV��a����&.���ڃ�F�'�������b���d��{i��,̶sƸ�����vӮ�4����u��lhK*Mk�M��s���'�9�a�Az��=��ݱ�ݣ�fJ�5�9�L�uV�i�	�P	x��]c��+D {,@ƯU@acP`Zo�����Q�QEN�TW3]v���Y��<�㪷no�F%�'�~{�>�kt��:�[�N�}N�^�y� �5V�eǘ�`�����F� b�"vhm	iV8˩Rߡ�OS-�����B��s���UG��5]vµ4��\�hB)y�g��Y������y���)�DV�=R ���F�� �d5(�����Etζ�$q�x[,^�-@�i5�r\;��ߪ���_H��Si��C�S��P`�S�^@?��e��We�0�@_���%K�d�mӘ�0���U��-	�K|s-�ޥ�q#�h�#cw(@���U����adS�B�b'w���:��͟o�k8E�b��
ĳų��s;`�������p|����@��#Ff:��dȸ���8o
#��_T�XUd]E�z�C+p�<�)���u�׽�-�3� ��n�U�ɡ}4z�r@�2c#h3����w�L�h�۞�,�(�/��B��}�#uypÉ�u�?V��Yn%�ԖS��p?םE4K�4���U��`�Y5;�o7�ALe9��EaG���m/�~Y�_=���ρ5�n &ۣ�������8�auu#�f*�XƩ�Ɇz/\͑�J�)�Ԯ}v�����jt��V4 ��i!�a�����
`Z1���`��f����4�k� ]�Q��z�ߐʃo��صA�����o-�}�N!č�N5 �����n.�%�k>����Ȋ��8��7�M�	��YC������	�jB^��	7��ܣO�Y��'�����<�OߞJ�����Y6��v�J��NI���a��-�����ɡE��h�/��5��O&)#����n���r��[�����:�g� )��g	�dݔ.suQ��q3ɹL./���j���+A�7�MLmC�q�k0GbfeQ����~�g��_���F���%��Ԛ�1�����Ԗ�Le�i�������`Q�^O�9Q)\V����,�Xy��~ù�©l ק���]0PW9eX�>��ec�-�~�f�7�C{�MW=֭�(JZ����R�ȅF�t L�B�����T���Ҕf�9a�����l��T��s=�n�	��{@����ʹšA��M��ؼ$�̝Y��P,}f8��HN*d$�&�aY�&.�O�]�b��j���V�y�����/�#0��q@w��a�TB��)�'����F�u.]���x���1
�3n4������1F��ҞNƷ|��iA�����H��q��R���_��`��������)9�7�LqXx���u4��U��o���,(��9���[b}�H���2���Q^�'9��b��k2�`����'C,���<-d�O�~��� ,�d���5ͳ,�c���pX���U�0��H��`��)Wsև8�a��a��U -���;�j��S�H��-M^�~��՞Q�y��D���@&2_�h;�:�Yc��~�(�*mŋ$�j�ùdh��(�Tɼ i}&`�o܄YʫDw�F�G�窜�Y@_��Gs��3��</�*)�;G�a���e���&*�����%(�;l�����ĥm� e�2�/>�j� �?����D	�v���O}�.eSM���r�%#�G�������"���Y��H6	��C�[�05�mO�����C�U�;�5��8Z��,K�'$߳O�tn�s�g�.mkh����A�^8:�1�6E����<�J,�k���"'ǩ/ݿ?1�
m��\elN(��އ��eq�1�L��y��Hs,_�ߊa8����,�N�@zh���)���y����w摮?n?�C�&GT�����Nʒ6i��֯�"� �r�jpc��|��@���[�G�̜��}z���̬����K=�=�mӆ,7����Y���,cFg�)�?/G��P{�h��JŜ ���+UB3�X|���*i�����͢|�΄e�u{��wG_
��������kvämH82�ɀ����_�, �����`�d@zq�<�X���M���������sg�]�R�2pz��g���^b�q@[����Pg���M��d;gx�0N�����8%,��ۊEC>�=��P0�i��eBӽ&��S��]1��4��h��x��h�	�ñ�b�WоV�]�[��-r{�u3}�ܫ&o�i�"/{$4xʜ3�����
rʅ[���0�J�Ћ�S0uoݘET�%���?�U`k	��ɒM����r��$��^Qy]K�M�&� 8^)*k��,:G��o�s��Մ��9.�Ӗz2���8GI���.Rk|���������Xd2�aB���p�����&����/3�Eg�vHٻA��ØI����h�� ׭�暋�r]ŌTF��s��ًoeN0�-���suį߀����q�.�Hb��bO��UӅ|y��'/��V<}��|���t t=֡0�����6�=��$=�����E�o<B��H;�	z���Јy���ed��|�H��*+�^���� S�m�B!yx����?r�ϣ�����
](ⱃJ!#un8t��S3��	����?�'�eTa���Y>3�������/�L��'�M\@�YD�m����3��z�j_��{P$���/$��>�¾�j\I"fK�E��rO�j����cs��|�����e��_�0�������~O���jP���	��Ձ��}�z��T�-��b�3P6o��C!��/Y�O�{��Կa�,@ց��+�Vt��s�����e+H��8Х�d������7���p>��v���}]�J�'h�<�(;l0�)Ou���ԏ���}�>$ݫ�9r4�G�Kɰ'ſ@"����o���B���C�n�Ҫ���)�Av�{����R�֔цИA�ƝO���GV;� >�u	t'��Z��W8g�Yqg�f4ޑ-;	D�`ߋ�n@{Z��p�0Q1à_���յ{��~��Z��3��Ĵ�!�ptЊ�w��
r��Z�D���t�{��Hp��p�(�����z�܊�,�H�gc�+�`?S��C�9���I��7gl�U�ڶ>����MC���>?ƈ�G��z���sg������=.�
A�3_wZ_Z&�]���E�)ͯ\�@ -k�;{����x��k��o����O�ցõj,�u��dr�0̵u���L��5��� H��B١⭎�PX���E��MZ8�� P��|�$}=ۊ���L�`ehᢅ��O��g��[|n�8�����ʛ�LT	|z�w�*�.����5�A����Pr|��G.�K'1� $
�
|s��%��+�1lFsٗp(�c\3���'}�`'M�J����cT��iQ�s�n���F�H|�B4u��n�8?���=��5���Bh���W��Y�BTץ=w���zv[��%��Q��V�ʒ�h��0&/B��h��=�7�	�;~B�N�-�-/�pPj��h��u�hUI�1�����9��],� ��N��_���c$Ĕ�`�l�+�f>��X�O���D�zg�@+mtӜ���(��շ,�Z�;����*��y�B�1OrC8���0y/�j�q�����=T!��n�I���A78����cq���_��#��������f��~i7ā�(�����f��9��f�Nv�ϲ��UH��G���C��'�v'zr�Y#OS�ͯyh�eݒ�_dJ�9�X/)kf���Oz3�gJ��@{ ,̣����#�k�%͍� �G�C�1O�Ùmԅ�,��u�㸮��M%_�&`�q��QF�`�7G�bXd%���-��3����6ʵ8�F�H��A�բ��]'�����u-q(��%$��،�0�_v�
36�"��?��͆��=�kxk*	�C�����^P��S��a9�Mww��.M#�������\߈��S�_�N�S١1ղ[����ƲqTF���6Й���� ��Y�Ifb��N�Ӭ܃��xTQy鵞�,~��
!rӎ�p�ϲ�A.9�U]牬�C6��f,�x�ҙ��w[-�ѝ>��c�!��[�?:8�OQ�:OY��x�Ʋ%8n�MN��]�I����2FlH�x�Ә�W;����Q�կ�R�i��Cqa�?����� 9P� �*l%D��ւyT�tvuY@��N�4�G� ��1�<fyK�=VW��!�j. �|z����`�j�bV&pR����/�'~��F�%7��<�����s�1�à��z�y�{��>�Y�.�O?r��A�ǯ�4��p��%3j/=�ߥ1�GqF�j�?^�l甶��"X���p�9��� t7���B`���夔���N�!!PU=��G/8k9�KΉ��w>�UZþ��3�4	\l�[T���@g�XS^��i/)�ݴ]Hᡯ�Gt`�T]�jG��$c�u��|	%ޔ3�/�,F,,U�8B8Ǫ�o��<����Y��,OK:'Z����q�n�<�g'�}��\��U%�;`�Ռ,cSo��.��z_�Od|�ӣg��s]���xbR�a�ɑ�(}�,b�h�HXo���\s�[�����,���A��r ��D�W���^o �(����󆀸�� r���4��Q�`��g	�Zq�q�ț��R����;8�>�����	���w�s\����y8�mZ�G�ݔh�W�ݐ]����!��°AAdZ/��ɢDK��6��FN[��3������c�O�5ׯ,��	��s�q��Kŀ����媢͚d��A?e�"w�v�B5
�y�l�E�G�) ��"�~��/e��^��u���
x�=�.��^�Nxʵ�D�T�s�q�΋�&zmW'���x��o��6�VG�F/��P|ʗ-?z)��Z�<lz��ʱ���������F{�c������ܪCШ�2��Pu�V?�hܦ��a�D�|c�O$��}��	)������|�'��x������Y6[�Lԡ2��P^~m���Ol�Ro"��aN��"D�Lq~�OvX�o~�#B`�O�~�����Ք��
rG�4�ݭ�N��%Vӎ�`1Z|�H��R�i	�.6�JܫA��J�\���[�=�}���e96�-�t�Y��Qf����l6}98�<��]|��"��v߹�O���9���g"�*;o�m��;ؒ����}i�\r�n�d�H�)�i^������>T�w�c8�Etd�����g���gb�e,С�љKO�:��yJ�8�%
��*x��{�ʷ+�7$�-�X(q^V�0����Q���̨����)mb�qȃ2B0Qҹ�KL��MFE�^�;�ʸp$������8k+1��4Xm��T7T+�xaa���"�y�3�3�5����A��H�T�k3Od���z����)_b�Ujq� ����53��4;��� ����1٬�
iP4á8��sW}y\��x|���²�@�f-�R�}}!�	�!�t(�&uU��2x�H8���OY���g��g-�J�#�*�>>�&�f�
������Aks�c�n e��~9�g���W��¿�5=�<�&ӕ��V��\�Z?�D0��8C9#�Ϯ��]LC��n�(�8s��g�6��<h�1�#��c5f!OOB`)m�ӷ�]r����fe���N�yl%(����n�`4���_�T�l�W�a-S���9K��z�E���|���K؂+�N&��S�W�}܀&��m7�3��1��[��~���E �j�Fz�æ�[�"b�f,��"�N,7��v�V�� R{8H���|M��<�P�6��r��.��X	/�k�D�f1H�567����}Z�:ձ�P���xt��4r��1��ȋ�d�鴢r��(�%�"W�a���_������c�+\Y>�
�[O�忹���\W,��N9��/	���ǃ�t]8'5���L�0��]x�yx���T!�'J�����+6��b�'�g�Y�ȝi�,�б$��@�n>���h >��qx#ѧ0�\X�aQ���%�4^�M��6���4*�ʨ��;NIҸ������$>�5��㟻&��I�m�"��,�ՙ���1p헡/� L��l���fK-y��W1�KhW>��~[שHݣn�^��u�H���}��70����i"xg#?���\웮uy0dkR�4� ����s�l3[���j-�k��^hg/�W��K� ��]��*q�����ѳ(F�*e�p ��`�T�H>{�=����j��d�L���9;�7?o����x��"�ܗqiL�\yYq	r�3LaS?���"���D��-yק��c	CD|�w��wbp��[�"-�_�r��`��|Nn�q,�5�XO������t
Z�Ej|�Ո["�f�n�R�� �Z�/Rϴ���^6H_��/�o�m#�6U:�}����GQ.P6ȿ�u,�Ȟ^ڻߟ��O���M5$�h��4���WcCq���	�NCy����c�"�Mʯ��np+,�S��ES3�����a�>�*'i�`x��;m���<)۔��3E���0)+3�>٧��6}�%������(�dxXfo ���Ϸ�x�﬒ȹyS0?��V?Y��lr㳍ߐ�!c���C�>,Q�����n�"9#L�������hU��� �cQ��O/[�����r�z�"s����f�MXj��ls�*R�$jm�ų���v$��t��m��CX����7>��'[�"�i���,8E8�"Hx�� h]�	^��|�G�W
�T���� zI�>���sOB���c�ZB�^�l�+1�b+إʁ�c�M_ujkyj����$5���ű�O�Ե��#�ρ��z��$��Ў^:���*z�~$r��!��j�56��TW�O�֑XQzi��� 7���1��o�;�����G?E�ǉ�mTY�(�����֖�.��ڡ�����C��S�J����IP��h&F4�����IV�� �%&�WoP�"�.;>3�L����T����y��`���BJ��P����f����\���w���!�BT�s���MG6&!W��? ��U��44^l��^���/KlV &��1a��2.�:^��K���a�0�?h�	�k3�x�4��6�=�L�r�����+�\��vGp�U�Kp�P2����3�	�H� p��Q����������w���k����/����݇�T��T�4�"��[y��� ��iѮB���sB�v&�gB��������N�Ԩ7`\V���PP���Ě�p�:�N�4Y�ԂHx����"�8�hY�e��n��n�Qc���_�����P�X�JN��;��w����N{�q!W�<C6K�&^��N�e(�i�i[�-2��KVy�k�w&a6f)�᳥v��K��� �\�
�}���=����w-�5ѿ� Cƿ�U6UBT�Q���j`hOP����jw�Up%z�v�%�A��&�6
u�n4y+h�ר�HDX�2����t������Ũ��"k�K�ۿ �V3��m�1o�7uq�-��xj��h��|�������*�Q,�~���]�s���gިl���K���k%%=�����ۓ~q%)�}��?�ߥ�.f�����(i3`��Z"~ ���~���K�@�	�k�@+�r|Aʤ�tq�Z�YT
���aG㆏K�ĸ;P��nI�pP��t��v>;)�OK)Ya�l�-�鼢����k�65�]�<G��xQi�:����\v�D[l���L�4l�%�[*�gqnX(g��|��?L���F�b��z�e��T�Amӓ��� -�3�	XE\�zDggI�.�6�
�wi���D��Nx�CR�J8��`܇'=6�W F��詈��z������?�vMh�L��.'aW#f2�j-[E�h���������X4�Y�U嘣���
�x _�+W��j?�!������^���A��j���j3�9{>�{&��_��
os-�Y)TFv��������.�~4�KRs�Rh;"�;�pr����K8�ʰ�R������ogU���P�>dբ!���#�+���5�@L�<�y�am6��Y�8a�D�ߞE�b����!ӮFJ�.�'�SN?<��)Au�܀���&���'�lw�����Ή\�c+��N=Fu�C/��0dDg�">SN�XĎvLn�o�$��ٮj8�F-�H1L�w[Kd��ߊ$�cw ��-�7��6��.$A�{"F��|'7�BK�w�^�����5�]��2(tm1�Y�	�잏÷)�ct�O"����Z��L�2�yPl�w�C�_�z�-%��gj{���2K��o�p�[����v9lS�&V�eZ�$�m�Z����^��> �9�~���w�4!RR��6��Bv��S
���}�J����=�5��M�ڈz`4·3���)T��T5�_I�c����苛�G���c3N��V�y�Zw�L�!�io6���O��D��=
��D��l~��I�t��]&�A��-l����Y�5F�Q��6��] Qj��1"_�Ɍ9�	���Hq�3e �e(LfT�?�?��I���-l������0$S'C.�����L;g�W_�G����:�4��@��N���@suX�t�, rT�7��J��Z��8jPE���eʐ�=���i}�����~�"�u��u��~�UP� �;2�����}���T��\�^�S�cJ�Z��nX�9=3�s�v*p�̝_���q4���2�����V��L��-��5r���zMn 9�I�	e��@���*���p������ǧ�v���۴�fsU�lI�M$�l�d`]zy��JJxͰabHR)!�AG"������-#}�%e��R�h�*�%�{�Z��ma����	\����
Dy�*�b��l,�r/6
:&+-�@&�*,���� X��I�p�RD�|(l�yeҡ*E�A*�!"ī�"L��P�������ί4&h9�d��?����aR(l}�>Mz9�1���B�Rn�+����� ��,Cy��1�%�c��֘LTy�-͏qgW�v���#��j��=�L%����^��Ԗ1�vH���ڊ�˭Ҿ�1(�{Jt䪚�}%�z񫺕@��Yr��O[���9��l���#a��� *� �/4Zs=�����i����l���x��wZc���"���]���C	��V��[xʝE�!5�ƻf��`k沁���O�)B�W��=�^�j� W�'��`��*^�1[�3v�Kl\.��Z-,�'�(�6R�險�EX|�,-�}��[�͠���y-L�t�/�0�>{���*��>�ƣnoE�	x"ﮫ����q�Z�������i�b���kn�T��Y��U�&]����(`���F퉭����U{�id���`AYx���y�������)�r������l=6�o&R^�?�����=S#n��挄lЕ7o���6ԏ2����y(u`�$�g
�w�;Lw��V'��9G�FrBv.��$�h�PH��O���vZ�=���]uO�{�z�
�<�����>U'Eukح�-��G�$o�akiqqO��2����0m���.}s�A�����(��5�ӏ�G�;��Q��L��5��8��2�t l`���
�d���"�|�>��I��8��w?�om�\���.p }Lߋ�9]�"��[aW���T���m��!��^�b�&M�b������$�ؤV��:�%�����Ws�f�ւt4F1����ŪM. �y��O6Z�^C����vI��֌Ҽ��J�4�q�M=䇰����/%����9�@��K�v� 2��ph\9�io��{��V	I����/�H��C��͍�	��k�	_�g~*f��-��@`5��{���\�Ќ*�w2)���}q���֝�D��,�O�ͷ�.j�EmQ*�����T^��	���f?l���e)�'�z�!kb1;|(C�H�w��ch�Aj���)�	�m��i�!��X���Nv�;3���	Z��rM�i��-���@v�$D�>�V�ZϟY����;=�4&���4?Gϖk�s>�#�V25B�r.��*>"�������uX��� "B) o�~����4�{��T"�� ō�rdК�z,�X�>�\$���̠����#�e2��@:�+y�k���]�Aj�%���Dz��sX�5~������^۬�s�X�!���F^�$M�h>{�t8D���G�H04iI�)��<{�3\z۽�\ޗ�<�եɅ���*�v�\;bٖgO�<�U����`H��[$\+������X�s�:�m:1��i$�c�������)ڶ�(	L!p5����gp;{Ty�ĘK�����kh�1^ย��m
CdU����N���iq��7yW���M(����;`;���L�ǢI��{��0�3� ����`���Iz<�>K9�@BD	�-��T����"N#�+��M�f�� ���$�o��RvB9n��E�:4'9��DG{��Kw0�����s�:$ی]L8���z����Rzn�B�-�C�����;�'A0#\[%�F�I�:�\S_�	Q�M���E�0����o��Yme�HŇ���}�� �/h�	
����TN�"D`F�3��U��+�א�<�`{|2��Itij�����^:�[M��y� ���3;�M����M�5�I��4[�A�-� �>A�`��D6�_z�]86Z��������%�6?��II�	h`N'K�vO���6�8��c�n�|��w���B��a�x����
�P嚊���bJJ?j��ﱵ�[&CW���0�������^�+?�U�_�Gd��9}��y��D8��"�����Rv4A^|�����Tũ�ڢO���R�{c����	�jOUa��n���F�t��1�C��1ғI���Ғ�3��┗�JI�S*h��6ߩ�����n��&�k�� "5�Űp#�܅w����OvR����s7s�5M���ʤN����8����/嶤�r��]�m�[��] <:����JD�m���n+h�T��o1uWA�O;a�@`5���]aaіZL��xJ�q9����y��z�?�E�|�%��n���:V�����9�%�yA�i_@��J�����X��?$Б��[�A�����64����J$��dk7�&O�;8 XFsw+���;����@�l���)A�n�+�<�]����j��'�Tv��W#U��2ȭ�YF�+.`�M�Ǚ΄J�딡�Rz>������k]�)��i\f�IJ�qK݁t�k��X�	�I�:�|�ų&@�����ޠ�Z\�#�9 J�ã��I������T��6<��Kb�o���E��.Ʀ�}l�)XXu�<��w�Ҿ]��ѻn��>��xҁ�%�%�r��Ξ]$e�/��n�$�ѣ���
Ѻ�PQJJJ�0F��
��B�a,�̀;h٦=K�����	N�y{�f��.W�dVn����[��
�|��-��ܞ��(/#�*�ƔE��%Ą�� ���H������2��V�u��r:�S$���{�$�#�:k���6�$ʫ �99XP.��V��AgG���ʔ�Ub�3O�X	B�V�c��iNQ4��3�f:ve;eqP�o:�����"�S`��e耩��?F���y��@�!͛q!ɦ��[z�tk.�r��PM��(�\�Q�n�J4��H�l>�،�=uޑs�[*+���j[�I�WZ�KZ��i��M0���N�j	i��>�_3�[]٬F
�0y����� )MZ���
�L�p`�Rt��g��ϳ4��q��/�=5�6%��VO���5���X�;<�#���v��{!�����B�I�Ɓ �-z}�� ?�DԬ4�8;0e���	�Չ�E�����p(����M�jo4#�obK���A��+��"������o�>����|��S�fOԄ��*��<�|~op�+-
_�I���匑�P�vj5��:W<�R����K�R�׍�sx��C�����C���@
�����?����,C�4rM�����6zDc i%��3��(C��g+ljj"���iq�����x��'�:|\�Ku�z$�e;c��F�uT��S����3�9�q��6��Wj����81��U��}���(�b�����Uق�Z��#�b"�hˍs���5f3E�e��V��CW�i�����b�z�j�Z�{���#ŉ�C���	GS�6�!���K��d�6<�aH�l��j\}1v�x�2@=��s���M������KjG�,I۶��#���Ҋq�fZ���`��QG(�����8ܖT�I�2����O4�U��1�������])$u�C�j�e��PJ��0DOYR�9J�~x3��=&t��|=٘�]��A��J�����	kMW��e��r�0]`�Z�r��Ǹ���T��ܥ2w�ay�Ve����䔿dE�ܤ)��I�6ވTywʢ������MF��&�vq{y����6�Vh*G�Z:���u%�b=�LA|�Jĕ9��A;EBEg#����h�8��Z�|F2���"5�Ϋ�C$JrG^��M�)،��ip��8oJ�p��	�N��lE�5�_��2�'�����rhV�W/����лG�@���ד��>@��E�7�,�_Z�U�l,T$|�H�M�ƧE��6� Ԛ���O�ѐor�^��]K��`�E�r��ҍ�ُ�Vj�#]3#
w��]�F�L]Hd}�>;-�������a|S��M?bk���]�G��
�xQ*$,� 9�,ph�/�p��)�@�S�A���Lw�8!_�	�cS.؈
W��W�B	s+�1�]y ̞��1b�x���<x�~d+��=���s�;rƀy�#��r��R�3쫲HP��߀djZ�������Q�E�1|S�/]Z�����Z���{�fZ-LU�#�G'*�)��=S�������F]d���X5Ga�$����L���F �Ʋ����&~�}�wC��Y��3c!b�i���􏾝�C��^=H���F��{��u���uI��=��OAb�e�;�]�%��)1�PE�W����K� !G8EV�W���oL��_w�Y�]�(�0�"b�<��&�E[�ų�/Z
axU�)C�-����\�������Z���~6�m`��+�vЪ�4�Ugqf���vCҎ)��bE?=���l�]��������1���f�ձK?��d�b���%����sa��g�0�_�1��dr�ĲlS]N��"#c���5d(��q�(g��=�[J:�.�w�f�����Ȓ(��TX�}3
�|�h9"|)�۾��fn>�添��=�V�����2`E���P�_�����
�:�Q?]����E�J;bt��d����R���-��$jS~�[:���tM�𸠖py/Tq�\��Icl.���}�N��C+y��DL⃚&Ҁ�ŧ;��B���0�e��K���O�p�-�����H����V�����39�2�#`k��v�c͍cd��k*m�*]&���;>Z��8���Qx��ؐ��s;�!�MΙ�c.A��R�K�b?��$�B����&B. &L7}	1���kS�Ī��`[j&��{�'b/���gaշ8���&Q��F��@���Wq�]V(y�7G���.�3uU�����umx7���gNHu���y%�y{�p���$�0�Q>�g�X=���m�3�A�A��[���"��˕���Zb㙽0�vy �!��.!�[�n#�4�]�|L�ۇ�{P[��@��k �v����;Y��4�y�ޠC�sǨ��Q�͵�g��fS)�4�j�Q& ��������u��[�jϐS�0�=wS­mW����큚&���;!��o1Q�R�����ir��3М���µ�+H�����a*���@��C�a��%����&��,֣9��
k
�Ae����ͥ��ux�g&>���D��Ax`��go[c԰;uT��7����7�����`lX��?CקE(� f�jt⫀�!|U����>R�(!Y�O�����1���~n�p�qV��u��V(#��FE:DWxUw��r�=^�gf�l8��O����qQP���I���i��U��Qy�蝠���Zb6�-n�Z�^Z8tG�����^l����
C}�R�z�Ю���.�8��Б1�'�d�4押�g6����3O\�}�6��e�ԗ�ۿG�a�ī-�S�f���E�l6 D8#d��4�\�������N���N����a�0�
�{�t���ڟZ�1'5ύ����萘����l_�n�r��4�#��m`}R�5.2�O�|	��B�W���b�{K]ݨ��<R�E�� �26�;��X���;E���D�>����Vȝ��ؖAx�;G4#���[��b�U��@�U��T��,@��k����D];S��FTJv|	$�"<o��;R#Ę�8��9Л�2����s���(�1�4$��S3U��M�h��>�ό#�9^�OTZ���0�Uym�s]�IF��00�sq�]]�`�,�"��,�
�S�`���)��>�GO����Pޮ�.v!�u`�.?cħ-%���H1�Pq�-�q1����MHgW��:ҿ�"��~~\�|{pk �ئ�*����=��J�v#2$o�l�2��!JH�y�_��m�<�Aln�hi,�ņexW[���vZ�5��)zN+P�G���n�������|l}i���'�CK��� ������K��k2})!.ֹdz�/̎<�H�#�e���o��H�I�k�s�/�:����(Z���~,��P�hȤ��w� �]�Q�{�;ǐݟQ4����U5C�O!"��_�5��~�NoԶ�Jx����OOk��o�yU4��CϥdF��y2�#�.n�9];碑�/1���|�y�$>���J,	���M�mP�L������m�Q��42��:�DR�`✴�Y�
dVK�b��	95K������iB�~{S�<;],٤kJ�F�!Z���������ɠ���A�ު:ٓE�;���o<:GT�)�"���\,`ͣ:Sv�}�>z�8;�`���	˟஡�`n��|F킼���E���e�{Ć6��W���
�W�pO&�)�j%�� x�� ;: vG�c�'�a%a�K�ꁥ�^0�/�j2ۻLYXp���Q�UjvS�%��9]ŋ�N6t��ISѥ=�6���{L~����-n�n/1�˧���d�I��:̴�d5��O@�!bGw�����^��p/�^)F{��������#&z��%�"&W켧�p�9ƫ.�ֺ�l$��8�:-D-����4���v��`-ŧ@�d�l,��&�HU�XY�4�._���R�C��R�>ϩ��[`E/�¬�[���S:��O�`<6�v-����F�#�ЁY���3�����g0Q�0x$)��}<��S�i�7�}�˙?u�c~O}_�盹Q�@� z<��Ǆ��gT9
���v���7m�
Ĺd�u)��4mm��4@���r���w�r�c����V���C��IE4�4-��d�D����N��m∜z��3.˕ɴp��v	�Z���\��h�"��	o���������@��ÑU9�����?^�<��+�V8#��#�ԋ u�4�_���b���#3tSƮl/I���)<��n�i�S������^6�H�^��t�.���_�NI��V�ovL^� �}��P[�4z�y�+  ��g�Hˈ-���r�v���q�j1@�Z�o�⫙{�ymW�q�GP�f��\�
 W�������S���bk��S���&���]r� �1�L����/����~g�������~��G,�ܡE�}�1rG.[�x*h���T9S��?AFL��YI��K����#h�)V����� ��Fm�S�3��5]�<��0�D���u4ͻ��Y��2i��S�G�c��evW|�:�CfZ�����S2�����S;�guA�VطJr��H��!�l���;ل`��P�T�G��~|�u���)��h�^H�۶)Tv
�4{RI�P�t��}:܌�(A������#V�Q*L��rx\*R���e���_^DA
���8�����2�2n�X���L�la�������)I�&�_��d}��ޫL�/ �l#�auUnb���).|���e�q�B�7�0�K�j\�A]�&{w�鉙<��O�Ҿ�P��N��x�3�\e|u'�	T6�k�:�����완Pu���V��ļg;U�*B��]�E����^��fU|��N�3�j@h�X\K��}և<T�7
4� -/�]�����+���]v�LHO��|��ZC�i�G�Aιo����'Vt����oFE���+;���cx�ۓnL�Є-_�yl�x
OC��қ̌�ֿ
@����ܦ#���} �ja2o�@�J�/��VG+����-M΅$���op���6�`�X�s����/.���.P�Ѥ�y��� ~�`S��^{O��QBT��[�%�Ặ#���N��D⼀7����O�߾��{<:ńoZ���dB���}tigdXk�K�j;���q�n��L&�}�8�N���7��1�vґ6c��v��\��+�ߓvk��]D����Z_Et��-8|F��pwv�+�b��Q��J6�x�f�I�r������1ދ���8?������Iq�����v��ڪ�)�Ὸ{�݀u1뙃͗��r@[��fe��F\�স��ӗ� ڟ�C��i�ﹿ��6�*��a��(�`�_%>;i磐�#jlA؟��m=[�yR1�H�e>q[7{DJ����#�E�vc��b1S�S���ͻs�@7���%�f��47fRݷ2|��v�F�[������\=�
�4�7�2����D�t�D"� %����WB:�-�(�n������tw�y�%���b������#�����0^��{N&�g�喍�A�ゅ���3} e�����o�֭��2ʻ��VÕ�����$s�pDM��������ѕ��'�C��n���{<a)��~���xO$�s$��e��C,��Zy����:at00��uI�qo���1�#n۲n%���e��v?�>���ۜI��C�������)"���~��!u��N����X�M���#��@��R,!»���#m�5�,x� ���1����:�ú��9j(~:����Os�_ݮx��@>��abv�q3�_ߏi�m��J����s��F+���1�Br*?��T�G�V���=�	�Gwƈi�E�����ܖ�0��s���+.���6)�r�H��z�/�XPR���\���~�H���3�U7d�\�V_�	�O��蜼4����bs^�o�0���Աs��u��. �)�u��&f%�hψ�t�XeO���Κd�c\�����y<�7A�4-_ͤ�z��7��|�(`���I$˯ڏ�s���EHXc�E�������������A�%Z������
d�X,�G�h��%	��U�D�Ո��_�i�K��M��m�c�b�RUzL���U��r�É�9�b��f����;
Zo�(��?z)spy���O6�����A�lE�>̃m]��P%0GL�)�x	�Τ�Q�rP���@L�1�5 d8pj��R�x��s�N�Q������}�f!��٨�����K^��B�2��`�)P�tb�_��6M0�]V�e$���K�]9B�\ۆ�'P͝'�U�>��}�֍��	�֗0 ��[��aby5��`N�;� �"S�w79�le�U�tt0/���F~���ұ���9�����ĳZ8��J�)�;�C4E� 3С���c��X��������O�=Q[uǸ�<xq�%�ˀ�:\&��Y�A�d�U��GhY�~" l�b�eف	g0�LD جP��k�Q|Ha�����At���.�ũ:.�bR`�z�-=n�Qi4K�혁؏^�0~�h�A�g����	U�l��<qt9�	�+'��O�e�Y��1��f��M�2����q4DJ-w��Fb�/�L��ec|0por�D�4Q^��6����e��wH%�'o���v��������E���(�F�3��e]� 5SZ>�ʫ;}E��=Ќ�d	�t�K5Q@Ut ���.��H~ x��I:փs�������g�A �J0;��i�;�p�A0P��dXю
���)�O�O�������UC��Q�]�'{���9��< ��ػ���H�[����SO�Ga�����l^h/NW�iS��q�9=f�K�>�#��*��,a�t>ζ;�+�g<ö��h�����{���6֢���I㨭ȶ2$�Q�%��Mv���O���o�\�'�gE���(T+f%Ǽ+ǃj���f�&&�S��e��}��j���!3���D�%�(�A?�4Z���><.�l1�%���|"��Ќn��aU��?_u=�!B6�0������ĬT��1�b�~�< �}4���j��(%������{�6��1���Ж�{HR~!9C�لB҃%}z��DC
�c�C��}��d����y���fO�uLk{z����GMH��i���Q�k��z�-K�O�opAiBkp����Y�I��%5�Y��?���M! ���y0m�c�.�Q�#8�� (�\��i��:�-a���o�73��}�^�jL[И������F�
%=�2cQ��� ⍊I+Ω�f&�R ��`�O���$lFN�bC
�����~�b�^8�@�P�ڥV#d
�`�DGlު��h"O��]���'\B��5J�9�𰕻-�L�?�h�|3��{��SX���W�ýo�p�ǰ�#��v.������r`x���{417|� ł����ţa�dU;�uX\�?W���G��(���?�YfE�E�P:�?W�"�8�?�Qc�+e(��yOR'���7��&��Z�_Nk�x�<N~ޔ�&�s`{ר;iu��fq��z񌺣w8q�A�pi�Y=n��o�X� ss���_�l�&�&2FF&�?$�p�b-�@R8l�H�!˟8g��?]�#�D�h��sp�9:ދaIn�L�w��p�m7f+k ���J��~ȓC�+TY ���?M����ʬM��h�ſ�SW�A����s�<O���~���x�Ʈd�U�6jP9�Cy��/�x�;�"r�����o^�����L��bx�������9=��`�Mx�E) t�/���YX�SZW}���tPx�{��&�����7�w�,T����`?M�]��ۻ�q��!(Z/�5�ٽ֑4.zJN*��4���H"]XAt옒x����~}I�V��L���\�T5��ǤT#;�۷'q�"��fBbʫ���8��+I�{�?I�� ّ5�;zni_ٍQ�"�T�?�����F���M+�C��y#�@���X=k�UȤg_9��Da�k͕��Ws6r�gjA�3����\[�n�`�n1�lR�D������[�\�zkB=%+W+НL�hpU�cҚb'��+����o�����0B����IK&p�~�mE����L�2S�0N��H���?�^���n����H^t��h��h[0�ْ�̮�Ġ+;��e�Y4�O�n�	��)�qz�]$���/.I���AH�*�l��ú�f^6��UU���&���E�t	�'��s�G�+��d��� /�	�^��N@�xHt�#7�Zt2�d;gモ�̃��!C���_H���S�lZO��-57�J��%��l>���������Ř^i���1�KƜ�B;ϻ�.�ԉ_�k��ע�|m���i+��}5��&F�|�]��kn�Lo���P)�ƌn]�u�q�	hrS�E]X�H�p�~*GB;�LW��J'�h�����*�Ryz�����/و�u([g{4�^;ɬb�ޭ���0��I���z�N{���
���ⶅ�Dn���_�������!��y���7 �%���,)	o�W��f����p͍OE������'�.�-ϭ(|�*�)>���|����2���Y����#�2Lжa�/nE��	��]g���gE4�DM�$U�6ZuӨ�M�:�~eh��
���#)fɽ2#0.vG�]������SY5��5�9%�zg�f!|���l"G/��١��3-�(�vn̷æ� ^m��-�*�Y�l!��7�~9*�����(�)�M*���F�����w�hX��M1�'�!^�3�j*~�ZL����`P����G	����O?��}�H%�8>vwڇ��KKD�u[��O���e#��+$D�I��ȼp��k�j����}S��=��UP��Hu����3�@17�ℜ#���^c@�¡��JT��C�/V{^�I���6��H�r ���'��z$�9��V��>R��D˸H��>��`0+���ԖR���G��)"h־�I	�f��o@]?�p���Ō�v ����ZO�)l"�Q���M\7�8bp�ە�*�3Jw����ʴT]=ٝ:z#(�,�c��0`�S�|�}�rLC�`*VB�����͐_��C���t��O1a�$�jW =����*����}a��g��So�T2���.�E=�fq���ش�.���P������1��>��Y�+�e΄W�"���`����;�E�y�Y�0�X�=�^d�).}�3��1�L3Jg:Gd�]e��$q�i5:/z�dr�"�u����̥�����,U�ڐ�n�,Cz_���53�Ak�*�0_�o�硓s�I�'Щ6/�ܡ�Ț'�2�����Y�4��L�1��a��6�Xt���6(�|H�?&�6W� ��P�9>RZ�تN}۠}<���e���v���p>�҆r���k�0��?Ƞ�t��D�l�`"Dͧ�N������Y����
:ה��y��q)̂ӷz��T���J'����(.���]�뿝�{�J:�Y�׮P�O���Q��94��  �p���Qh��G&Q3}�������'��!� �>Ba?���S��f�*T$��R�����8�"�u��6��2!Dy]E���C�ہ+�v�
Zȳ�e���:.��kq�b����k��\$�k����cNc,Wb�Ð2[��EAYd�q�����V�@�ʽ�Z�%�VQ{y>J3�K͎~(06볆�N��D��ȲE�t85Q����xx���Q:\�y��!cd�6m�P���P�M�U��kq��/]���b[2������0c$F���$���f/Xܐ���	$&���F#`e0?�	a�,��qV���g&
'��C����a�>2%Q"�Rv������H���y�i��?8��É�-�86wq��3R2a��%A�Y�d�wo�k�M��ܑ�����^����|�ֵe%|���]"��K��ۨɇa�"VN�O�^z�݀M�/�h��ȁ�f�H�|bzE�9�n# d�}58���:	���d�r� �k�����Z���\�S����	��I�I��+R���N�v)����������1���e�!V8֏&������U;j�r��#���iZ瑅Z,~����G��YhsW�ϋ��˴���5��E_�Gð>�Q�w��2;:�s��=��W��xVnk�ՠ*JL1�qAq]y�-`��c���@�;����(xY�� [�'h�b�O;���d�a1�;�xf ϋW�,�JN'�@�� ��j���2��	XyH��֦���֋����43F�3�^�fRN0Og� ��Q��7Ğ�߫I:ݲ�D3�3����'[[���^R�A�s�N��frUk���v��ؐ���C[����g����x��(g2��<h�h6An!�J���P�����R�(*�e\ʁ�X���s.�z����H�����H:����-������r��(Y�@��:�:ÿ�\`�ɒ�!�?�=��������)�_)SN�j��� ��>�������r��s���Y\q�:���s�΄�tʷ�Np�G�C P�����
7j���8���{��F��[b��	�c�=��M]��:l`r&��B Qi� 
�j�8��Սr�,B�E+�An�1Wy�Ԫ?`�RD^��-�6�=`����6��P�#ʋl~��ݣ����]=���1�<PϷv���ƪ��r�ʵ*�X{&��q��d�
����j��a
��t�h�
Rb�l^W��D���P�j:BMokv?E��`@&:� �@p�?��~�~�u��ʚ���f�B��U�y%/�4�5������X1QĜ��w����w ���ḠG߽���W�I&;	����97H�p�vy���-���h����KX43g����,�U�AX�_�f�iCɰ�D��@�7a%�..1H�*�W�M*��;<Y�B�*	I��ߜFf���o:�z������&��<�7X%��R��3�K����RS�.V�,q,~2\X�'��p@�����T���c~(�`\h�D!��(Y{1�c�jB�c4�^W@~TG\��*`�p��eyB:Q|!��1+���z�1��5&m̲+�7K�i�8u>�l�֑͐Nt�r�)'t42ղzb �!��"L�A��X�=���GC�K����̖a3��j�H,@{�W8p!K�8�H�g�\��~\ڡ��������7P/�D�;��N�U`N<��
�XM�o��%h�jỶ��W�NFoa�d����NfgԬ;��C7�T$�����urE��TH�Ͻr�6wd~QȐ�^��<�s��
�>4X��Q��9��^�~����}����T��qu���_��B i=�>�y���p�(`�Y��O�3�Cw��3s�����~��P���F�!P���ӝkG��~�5|���o���&�A���JG��uC���7�>�Y���I.��37�O�u�N�o�
��,q�2�h�����X�f���^' ��\~)vp�)@D�J+���Y�[
g�?l4�م
�O��iL��T��/�O}��g��Pf�h-��D��#V�8��qh�U���*}�����D��,�^!SX� �l�鉺�j$u57PܨI��Հ���d�ˤ��e�.�
Ԛw=μ
"��i!C=7�]��\�O��1���
���`���Ϊ{��ʟ����Paߏ/B�4��ʺ��Iȿ`ch"z��R#�H`*��JJ��w0=v�Ә1�{���<(���ݴ� ��c�H9���"My�����'r�^Ffh�<�}�����e�5Y�M��=��!���_&�)pV�? �o�vHU���O7偨�ц5O���6�^pj1����5�j�{�8p��6]Z3�{D���.����zZ�n�ưż]����=z)�u��,ܓrj�z��6q�s�d�NH�Q�4��8,�a��{Ö�	]z�kM'n@���f��� ����D|u|�Q� Juy��.����ӳw�+9BAJ\d���sK�A&	N�N����� ?�dN�w8̏�����4��:�`X�΀ɐ�d�;���j��38kC�y�J�>i���0�\�I��c�h��:����=�}8�f��a9�'�fw�-�ok.!�'�4d����Ф�5G�����f�W��Η�
9�ۜX�~z��\5^vBյ��Z��~�"�� ���p�ǩ������?�B}q�@�&��k̰(��/`��{�$�I$���5_5:I�%|7�t���z"J���4�Tv{қ�1�����v�^ޟ��؍�©"�%a�x*�4�b-{|���*�,Y�#-�K����8�KA��*�$,�N	����^Y�6~P��`����J�J�:$	)&�u���R��4�S�ɤ��� ��UN%/��7/��rx�]T����I��l��^���F��>��k	�y+C_���]V�!��0ٷ�;�qZ!��Ȳ|B,�̪�=�8�hZ/~�r�j��� ��y��>>��i߱���W��]��4��9�2��}}	�x��/:���!�TL��:9�Ω=�>Q��/��1OS��O�����{	'4��[�� '������BְF�hTF�GA�� 4?���ҳ��2�2���-w~�=`$������`J�� ��m #��>�_����t]�V"^�.���T�[C�2��J��]A��,�m]�����?��k�� 7��\���R�ᷚ����X���I
��*GYtZ�ecntO�m�=p8Q���dqV�˅� &�	�
RHư��nݠ����]�Kb��G~��i:�(�b�=��J?��s�É�W�x�R.v%�ʄdJ+� �a�޼Z�5����"|Y��,����	DNS�:�P��v�R������n8�o02i�Y1<_z��ց�F��ҀfQrl����xh�~?�%İJ�t��i�/�t������ך���1�g�A�v�6M��j7�%��]b���o�z(/����͵�+̹��c��(�E�U�(�U���h�L7 OD�wk�g0N_]H;O���p�4��6����'Kl��[&�xQ�U�L����p�*�qs������b�Y��2A��'�Y��6Kv�7���u�ۥ��SoKސ��U��Ȥ�5�=�W�=Y�s�&#�K�ƯL���R���+��wY�u�^�_�
p7Š�7��͙%� WnY���I�b*��⮭�|�#b@A/���F��� T����S�����]t�9��p�$/\�$H���&�6z���I?�w���S܀Ǘ�^�S�I��aG�f`^|����H^�0/�9�P�!�a�<z���<�zwu��<�L�)���QT�Cug�{��Z&�[`M�qf6@�YA	����,�B�V᎕͜���.6���oz��ӿ�0�U�c7��MÜ�e͘���	"SYE����*E�$�M"Ul�&���򨫤�\��g����r��G��r�+C�Z]6zB�Eۄ�.�I�L�A���t�d_�L�:�'G��꾙�t*� ]\��n���e(�8E2S�n�`��ikPћ��:��(���c4)ìnd�یg.{�v,=�(6�hy���W^ϧ�<�[�����/�*�ס�O�s�ꢲ:iۆ�A6:9�ኛ��j�c�����m��V� ��a
���}�@'����sSTK�X�}����!k�D�{��u|��O#��L�����(cn3|�b֜��T������C)X��b�g��:U���"�:����ԩ��d��k��pi=����p�t� � ̻��t����YB~�\\�l�6\dZ.� ���˰��t66���ْJM���P	�����6�O�Vbi<�p��9�ڦ��D�Zj��V1�_��[��O=6�k��-c���"�,S���-��X=�7�KK�[rӅ2D
��4٣�'(��9�fo��.\ۇ'U�V`�e�]�Ѯ9�yw�Ö���
�$�@2P�clf�)�Х:.�Z��L����繳��~��r���^`���־,'oӾq�+�y�L������ }��|�9�hg~�W�>E՗"����9�qx�A��Ff���V�W90m��k�h�n�~!��/	�����@�O��/��~���-5��j�p�=�amH��������;�?t��~����E$vb��DR��A��0[�&�m�tV��`P'dd_���-5�BGasX����wWN��j��3�CݭO����@��1$�e�s�C���?;����4]�(
�ԫ����dﬃ��E�i���	6��f��=�ϔ�C;X�̛�B��m�����t�#��T�	�-��rd�c@��w����){�Y0=$H����
!m��5�_z����w�������fRv�.M�)^�IH��	�|1�s��hz����Ě�3gO{�(r�]���0�Ŝ�q�k�P�G���}��9#ӥ����}t����>4/��&n��OT�4��q�|U���	�22��b�S��S~��Ѝ���F7Z�G�-S�S �j�sZ%s���[�QGY���!�8ųD��)�Rn0{D>N5�\&	�ƞ!�f�"�p��{F�6޵����}
@����j�R��J�8������U4���y١Q��w�sP��1Ma���+��������-3��"#a��U�����%��$%�Ut}�]j�	# r��D�Q��xv_�8�K-��*q�������P\3^6�KZr�c�����܅㶩�gl)S�  �Z�holV�5F�v�ŷ�8R�����`'�o%	� ���&d����k��ZR�5|���j�]v��v𠼸�ۖ
��ib��T�X(���.�'�Si��(�Z�����k�t,"i�N�Ԗc����H�n�?��G��ч��M����D�6o��[�u@+�*����k�MɌ�N�-J���q�4Z8_�D�}2���6b�(>��&�s��*$��	��C
�gW����I+��y��Y@���i��}��Qi�s��}GS��.-Ys��jt�Y�& �Č�m)e�$�L�Z# >���U��h����VY#�	�h��8l��WsIC�Pa�� ,��&�3gfȝ �"�vś�nJl���镵iV�ȭAF�r)ge��lJ,Q�dG��K�
��r��/���-25U��埱F�>m��*�Ӏw��}�MC1A���)�M��Xnq�d�����v$�*,��wh��7p߀O$�g���k:�Ŭ#�]�:^`��j��ħ���&!���F�b�pv-���"O^��snu��m��ܳ��P�FJ���j���e�,6^*�p���#)t�)���0���Y�P�c���yG9F8����d��N���;5/�+��(���󌇐�(�Y�L���|
�Y�}�3i�{�Z~���S�0�����U�<u���B>i�1����7�e8�Б���*/}?��{ XmT�>q4S��Qs�2.]�=��~M�s��m�)�j�Uc|e=|�xY=�^XW���� DIQ�S.ɂ��_�
WM5������{��t~�G�r��r��P�j2,u��&f`Z<�9}Ay(oX���g��������V,Y hS/�Y:��0e�4e��>kZR�����9~1R��u�B޳�)�qTg�u'#_��ܟ�݋֒��9R?�AS�1o��Hʅ��QG=A��q0���h�_H��\�Ƹ@N�9>e��S4��u�A���ن����}�Qe�-�k��A5�X�{��`���g���[��e4(�-�����񨓿7�+;$5:TC�@u	�2@���kr���s�gh'�����۩9��DgMQuʺ��gM�h1_���z	|�z��P��,��v��ֈ㆖K���D������*��9`�z����/�M���g�^��OpE(Z�%H���[��J��������H_�$\&D���6����{-��_�V��n�K!�z���⑜ͨ7-l;z��zq�b�kO���!��W�
��H�����#6������E�D]5o5%��UJ�巇���VR9����u�k!>�9����Q{6xK	-�+��*�@��Zm��݌"�	��*�Tkmi��l������E�5�.Ӣ��6h-(�V����廴���}A�k1�`I%[�I��%�^$�#��4���JJ��2�Z�mOR�C�	����ȣVYu�qf�����jU3�c|6^d�*s���D:�	�>um;��컰�g����C�h�x�Qȵ�Q�M��MB�bx�]�n�b_�x�8��?,��d�+v��:��h`����¢/���d�AO����kfL���X�VC=٥���;���7��Ϲ�e\X)����HjPc�v��0�>ƞ2_��9�
����Q�U
�t�����!���<F������0��-�˘���ŉO:i�L-�]�b#��ؔ��QM9�Ek[�/~6T"���.�� �蝍�.ߗ�a����.�������u�%x��k�j"�j�a09���FIy���Ki4vEt?C�t�DA�3hܤ�h���X��\f빰��{�R8�y�;BՏd�~|��\DQȲ8
��/ 1�D��#��@�^��xM���I�$���''��u:���89V�P����>F}�^t�O��
�éUH᫼��hG#�J*5�9��f0C�'�U=�k��5�{A�%�ջZ�gɉz5D�����0�Q�*�k���� n��Y����r
�z�/�N��8��� T�4a�e�m������R l�y��y}�MF7��(��,nHb_%b���/�OD�	NXM{$����7wr1�;Кw"�c�j�W�zՋ�E�~Wp�_��#XP����jZ^�V�Jp�n��b5-�>r�/I@Uf��b�	��2m}+A�64�>�'O�&��0�=�9i�ٯ�ZEY��vZ��U��K照aQXaOvדvf�B>��k�^�|E�G.瀠��`k>���X�]���_*���8�������قo�Bvf�Λ���TUb��&./W�d,a�=�E��R�}�.�JW<�S��(����m�[��*} M�N&��Ti�!���0�Q�7p��wo�g�N[a�\[�Kâ�z[ �����X�Uv��Z����l��۲h ��?����c2�q'b���p^���G�L���$aׅ�� �|	t y{,^� ��x���r��NO��������#�N4�h�����!���p�ʀ�u� b4/�G��ù��g �s�'5 Lg�9P6��k��,A[$��m�)��*���j�H"�݈EJc�H�vZ�������[ږΐ�8�>mt�彾+�s��xb�ܯr�w1�j�_ρY;�wQ�R-l��~p��KQ0@������c$' p�-��Br5W�ƿ�~�3�mlĆjVۛ8��]!�Ux�L0�I�q�_Zȓ?k��*�s���lW:�A�3��^�m����������B�<cӊDAdo9�粤���B��#MSڬ35O���I�<�==Fne��ţ�)���X�ڢ��S�o�6�̍H��v��y�T���4�P��3�r��z���Md����O^�m�휌Q�l�.�zM�oƥ��5 �6�t�#���CL6px�&��s��¡ue�����7&
��2�z������Y���Æ��ppx��d=�������M�Ѕ�?�o��F78�s��(Y�0vD�����D[1� Z�R1�W����D2L
���|l�:�5�5�\	!</�ѠVZ:@N��8[L�C.J͇���y�'�:w��&�B��yIϕ� B:@�����m%��ʁSXTBu,�h�D��+�rI�3��&��	G|?��Rze�Y_�l����+^&�Ϡ�w��I{�`E'?Ġ��v��,~zC��p�� �e{�\.���Ϡܮ����콐�m��K��%���ϰp�bp��nn_�3�巉�0i�~j������7ۛsW����\�&�������2q�X���NK<B��q�UY��F�/;�a���?'��oL����FJ�
eb�@�Xvd��E�v���*��0ݺ��O7��,qw��K4���Y������0��S�. �&]�/W��S��U�Vp����~���窟�����|a
�^�5*����~f�@}B+#������q��]�i25lub[�s�^��DEbeZS��w��Bd����E��D��rj[k[�g{�H1zy%#:�N�҈(���a�h�S3u��7u�t{n��m�&2�H������B��Aa�@��ڲ!���I	jܘ>{��|h�=X썄<�qYʅ���P�[׶D;�Ș�nBG�(��Kb��[�Q���B9g��[�Ws;�۬O k�A)�L�?� md-`��.���>�dS���ii�I"f8����h�l��-��!V�'H�ìQ�x|$����j�)�+�z|x��|����0�~:�St�\�̑��J�ft����C}h�r��^��˲=P���v>#a��*R��:L�}c������iSf�i��~�:;�eZ�,��̂�����Di(��#���Ï9!���$Q�	H�������x�����rg��*'3:����o����#	��'�q�r���F7���f٭�ӡu�<�n��k�ǧ��"��I$B�;*�뗉J�=-��P�� �'�G��t���ۈ� Y|��	.B?^������
䫙�ȦY9�G��"��~ C;�?P��}Z�_��'�G6}��}�:Bq�AÌ��dԻ�Hф/��)p��� �ls�С3�~�8V�
�?�w�I�� t�W"����P�q�9��� 	���m�7-G\}_�g��,Ϊ��xt��w�[�M�nEDv�bM]�2�����oT���s��Vڳ�%s�y��ඛ�o�y����`9�o?��`���
��gDf�A1 4�U��=��Z��y��Y�OoV����N�hcbhm1����mMn�0��@�����ca��|Q��	�aĉ�6���W5|5gq��R�a5׎���6�h8Ni��� ����@��l��@�ꔇ�V'SZBKWw0F!��������o��B���%���{�پ#5Xwo �"��f�yfFo#��^�|��r�5L�\��/�ζ� mP� ��U�������6�D7m��$�e�^��u��Vw������U��_���z=C<iK�;o���E�&?U�o=4L�O�+G�.ЉX�zt���>6ċ���Љ|}T���N��i(!(^ �>A=_�%92ҁmm�T�*m�C`��7hX�Z��f��Y���t~�\o�^�������km������bŖ(��*�e�%�N&��ː#��.���c,�����S����XX.�7��y"�����/�V�/� �ď"���p��JBњW�Y�|B���sf�h�@�c/��5V6fBԯ�H���u��˰�᪪��kO�1�!�:�G
_|�Rદh�b�8�0�_��oXV��D�N$�.�����|~�{��e�A����{��ِFaF�/ϜxԴl���ËDa�5o�0��������D��]�&�㼙\a�6�dv�����e�k��H5"ڞ"������8.-tv�	��2��m�����Ib=�D��xX��H���c�+�9՛5�%9�9�m�耦#��w�!���0˞��<�|g���ҟ�:�j����T�guH+1�f��p1K��1��aI�3$�uS��Ͼ�]����+Wīin�\���R qIӃ�`���0N�F8̈vhM���wk��ܕҟ|�L٘�z��5Hq�ȴ&�o��T� 5����c%3F�T��u�$�+�� Ep5�ٶX�E����ugZү�O����M��o������<�Ά��V3��|��@P�Y����D. ���m�`*������~��H�qDC����l	Ǟ��$�~8IY�\��ȜQ��,�c�-�!�Whm�A���X��^w�w7��=��M��!:0;Gx��������?�v%���M' A���[�P�����~ �0�ώ�5k�k�X�6�Ϸn���Ϧ���o��c�;����7�NK[�c#�E����J۠���:F�a~������^�+�܏�v��;�|<�阿t$�e�7Hâ�*<U�D��;�Hz��"~�Y:�U>�Mz48���W��"O���	��1����uFޑ���/A3�6�.M� ��!-h��~fhB���a�'��]�ں�V��GQ���b�h��5;��D��$�7x o$)R���{p��CVB�Y��dW-ܥ�(�Q�c8�s���AT�NL��G�Í%��S�8�9��Z�v�	�=�F ����J��+�ZE��B�XRS���K}�a˩�XR%1�����.�,���ZQH�9a�AjΧ���Ys�����D������
���� .�0�Iu�Q�/6?.��t�O��!J(K��A��x4��Fg�{
��k{b�^��ϻ�r���7I ��mC��Oe��9��-��􈒖J:��O�t����a;�<0�����"П�1F�>e�lYr��\S�>A�-5�z�`�����DG��B�T� /E�zU��r��Z�CĻ� ]��"E������C��%F��`���
���N��O3�V
�7ڄ
o5{��62-�T�7П�»����=�hKqb֘k�b�x��_�ƸBQ�\��n��mI��GB)�YYm7ȱy��oR��p����i[�ueU��x���P��Z�e1��G�yt1��
v�R���Eܵ9�7��X��A��M}4��s
��U�\�����x����a�/aod��m�����P�VJ�V�Ӥ+c�+�_���O֊B�HA^�C�,F������9�t97���E�_s'�S��[����۷�JJ\>q�x�E�B��;��ԕ�ȡ�2��Q�M��|�����XtaԀއ6�ȍ���z�'�4[wWk.��V]%�#`<���\�UwP�C��PWd�Z�u�V�j�=>1Qt\�B�\��X��R�(�m󮵂(����y3S��o��3(��t<��B��,eÎ
Ym�ɹ�Pw�T ���~���~O5ͬ��rg	#U��)����ݻZNں]|��gi�m�������eG�NU-���O�|w%�%�,%����tS�$�h���m?���t瑁�IЦ�c��:b��n�籘n�af�D����f���m��C�D2��c�2[lT�S$<�S��G��Ij�� K�����Ł��v�Gu�'�i��}b��g<�~KG)�$���)&��I!pL5��a�׼� 芟��e-ib�l�i� 7������F�S�!"�jz4��e��$e�^y*#�ڿ�{ &ssf�.y��	*�1����
I�z�m�d�;��v/��<���-T��D�e�� m*xFa��{ef��`�쩢>$"�\�RgF/�z����Em֫�*�Q���w!L�%B=_\n�"(��R�V��̋��<����;b�U�NH/��ݓ@It`��W���"�D��.�R@� +����L��z���?��Ѯ��3��:'=��ҰY�<�_�.x�D��:�B7�Ƀy�Ig|�ͅ75��RI���Yo�;p�g�9�<�o�M:�NP2�����C�>-�ݭ�f��<��������U����G���R�����'y�������(��<Y� ���+�1� ��ȣ]�d���$y����4}6sΌ�}537ʞ�+8�Y���Y�Mx��~�!&i�+J2��V�ADd���hGL�@Pw��nN�#�GT�.�X���,�G�R��5��i��@4�Y�S�`�Q_�	�%%Ȗ��Y�Kd���J�Rcә�����٦̄<C�`�ȣ��z	��Am jf�kZi�qQ�m��X@���i=�Kyr^�}*�VrT܈�M�Qw�I[�0~N:��ȟ�#�J�7q28kd�F�ڷ�б_�~����_�iO勸�Z� ��Ȫy�i�[7�$`u�y����! !��h�z�|t�����޿}��i1���k��lu-�7΅h�2�V���%2����f��R���b	�~b�Ͱl�{}��u��a�v�qHҡ,ِ�3�4�B�M����G��G�
�E��
��49-7v�s�\Kp���������Q��7�h�jux�v�3��)k"L���wX0PD�^T��5KZ��'a+���B$�i�����i�W��;u͉����F=a�Jm�`�)���~�yN	vO���۔bjb�S��;�����eX7\��d�Q��%T���4���H#��Ԫ>��<�IwG8�4�+���_�S.��~�E�ͮaQ";K�W� �.fe�^.�8��Tf���Q��R�U�8^�a���sD���u��M����(P~A�CЙr�ž��$%NƁxN��?�}-�-0�/�ܖ�f0;���L�N /�_�i��o��ْ\�t�]��&�@y�������`�Ç!kC3��������t�uj�n�Ȟa�Y����s�#�,���\��
۝��j��w�f0[s#��MآXoaG��7����D<-{��u��	|I�V��e�RȈ�*'��5��}-{��g��7�y<���{|�O}-��J��X��>��l�Bh�A�Ĩ���"�]��ny�Zz�O���>L�|%���N�۫�HB�e�s� �4y۪��zsժ(d� ��+��m�S���][�����a��1�Cȏvh^O0�XT�m ���q_���X��z���$wW@�ߋ�}�Br�"�����tY# ����)@�XT1�����2����Ř6|"=��d�/U\�����r&|M��2 `��[
+A���$S ��D-EMD�J=����G5�*��+��NӪ���0�K��|綽�?Xa�Q��6��P�tQ��ƥ��հ�:In�>: m �3ۥ-z�,�MGDU�h�O'�0�M%l"�K�LNP���l*;���7�i-�1=.�/Jd�6�U�2s7g���BW��!G�%	!�?�jPlJM�8Y��{Xc���a7��������G'�tD�>�f������Fd�J?Ka�!	E�KCa�skY=�+��+�J��;j��M$�9RY|T���ʂ�0�w�&�)��;�O��w���8aԖ/����aI�FbsdM�(}��N���[�b�i��0���N�~O[x��v�������a#R����V�b��}Y���.TXR����9�6�qeyo[�@&"y"c_��.����8��FD�ФZhT	��v	�S�vF�CH�pX���w �)S�6�
�5��t��^�C���y��D��nJt��]R�$v��V=�>�׆pz��}���IN�:�5�=]:��4h��
ׅc�����S�@���yH�D�:��xr��R�yU�r(؜�Sb�r�h*��M(=�*����W��5-�:Z���4p�WU*G�:U�qoT0��P�[,�,ay��ǹ<��^6':7(��f�k+-Ҁ�%���㲎��Z��-�q΃V��;#�V`�;�͐��6������˔�(Ng�t�m��I���v+�֊��[��=�&f����R��	���U� l���+Q���(�Π,R�{U\FG�	�/h4? �y;��F.�ڌ���}N��=-��Qw$y�@�8��
]�����
�	L�ג�}�;�~�'�{h�YC {>��u&+�%w������B��
�rJ(D�Ku����5r�wP�+�
U���� j.���u�Ш�ZGw�HERB��)[u�hV���O~u��l4z=�縸4)5����9O+4�|�@�M^۽��Zw>qL��״�+�7�7/��)}
L��$_�i%����f*m?�BS�y���
2p+k��
�9�
�7I�d~ɫ�>�P+"������5/l�B�#&��K�|�HWt:�/�Ќ��&�$
:��t�_��#e������w�� 1Bs-͞�i2x}(d}��7���[�E�*���?����{Ah���~�Z�a[�O����Nu�09㴔+U��tY	M��5Y*�n��/Vݠ�ɏ�6i ���k&�X�ʕ�]��I,d�(��5BI>D�i�,{)�O�� ������|����x�Fˌ��9�\�"u �����AwD�2�����"dc�<	Q�� (}��p��}8�8��Yo�@�<hSaĮ�.�J��F�k�������cG6�d���r���u��J-;�9s밻aSH��`D�|C��\d��g���m���JO���ڢ7k�J������!���ؚ}Bj�C�Msi>���v�˥]m��2� +�9��S�����h�rc�����a%�g�W;01c��lE3�՘.<�ۏ�t*!#,.���&5�'NK�<�@[[9i�u���О�������\~���!�i���T���7��T����H��0�ĩ:���v��p��+`��&����ή=���+�?A�y�9�`lM�2�V�dnhe�4]���®�/RG[�y{���-8J�8|j�S2l�G�`N�>N�;PMɀ��:ˤA�m��Ns@��1���)t�TO�Da���%C�*u����ÞJq�,[b%�w��
n9��)PiY��g�6k�T���ä�I�$>�m�5R��.���bb)��?�]�2��~����L��(:w�
� �g~�4�n �լ�E��YXۑ���(���h�VP�7�@/H1�o��.bk��3��X�钝��0����W�#lҧ�5�[�E��`!��Z��ܽ������>�JwA��HE�.�'PO��`)Ԡ,x���M��ɂy��y�����-г����~y���@.o�C�ÀO"A�Y�p���z��if�L �V"��:a�Zc�4JV!VQ�5`��;#{�bW/մ�^���X�?�%Ε-�9�i�7��f�t�b��Z1jN�!rV��l�1\�*��<6]��a�<��a��{i��f?�j���1�:�9O�/jo)��JH��r���������R��J*a%�u}R�N��ټ-:Z��q��!�� |�9?4��ھ]��M%���Mb s��搮�|����b�p ��A_�n���V�X)�R:%�i��`�����mܡ:�(T��u�{�^� o�g��q�*n���R�n�i뗳�7�^,qkb�S�V�h�{x�c�^��;kG�Vuɮm�xF�����C��"y��y}�{)�MT]��+��wzd1������0m�0t{aكǀ�֝�Lz��lf1�>�"��>�i��k�Wot�PF��ݐ�(��a��@���W���>����E��ܘH0DIwi+۟��c+m��Ż!M���iѹ�]V�����܉_2��V��Vh⒩�H�$�s�.�ʊQ�T'UC�ޔ�F6�f5�A!���vB���t�M�#�r�av�'/,$�L3��V%U�<���>��	�zȢ&��m���з;�tA�}��d޶��E�w��s$�̞�,��O3�=�����Q�A�	���d�E�pU�e&2���ǻw��u��v-�����P�`$��@�^�m�&+S�|�S�셃�Q����3l�&&p��#a�F�ȇ_��V`DA��YVݷ?O��<A~����<�߹�S7�H!�2C��Le����6�\�#ԭ�8���7ʱǹl���\����,M�dQ��(�\�֫�Z�yK?��u.#��������L���;[҆�vh�ԩW%���	p^N�(��n��v{�?/>֊�}r��$�>�]�*�I�
Ój�V�X�%M��YD�Vs낻1w��L^(���gv=�(�v����u.k��)�vXR�����K2e�%1�2�k��U�����g���*2I��r�''���E1�cՑ){C)Լ$�(���ޤ*W�Ń]��s���n�md ���Й� �s��w$����)Q�Z�x�UV���k�A���VT����n!ô}�NF�+������Q�eߟ#�������_��{�{��\rFs�X��?V��=;#̓�/�O��xY��9��l�Ē;�p8��'���\=L#���p.'�'�u5�](
���������u�	��A�"^�4�ؿ��ik
T���u��&8�="xh��ә���l-:e�F{U�X��u�W��W���f�X���ɵ�9�� !���&4�FD>%��vY>M��Z����A�B N�Ð��wDP�n�؈�6pث�>�w����,���.�
��9ԕZ��x�T�����^m]��L�ƩT~uG��>o讇���"��3)���8�����ߖ�U���r�����'p{�ٰz�#��icGHdt�����h���[�}��]�1a)�m�9NWR�Z�E��UR��.f�����x��\R�i�'��^p(c�n�$�37�zz��E65퇯:K�bf�#z�>�F �`vn �~��{ɠ3�J��6�8r�?�uQ�.o���o��5��
��vR]�tB�Y)3z3{��+b;Iɨ��5u.�Z�t�}�.	�)?X{W�Re;F���ط%CH�a�j��C��5d�D��!��{�}4����Z']��L�W��i��~���&�)yҪ��CmD��T^9�{��
!�%��Α�VW��nȾ��eK%�"l�_�X^+Ɓp��4���-�WTXRp�y۽�q����
7����_���:8=��D�r
1�V�7�|�QQ�ǚmƠ#�1?y����y�ΕOf0���N���O-�@-<
A����V�ȿ����|@�Z��+y�\�1����he���"��7��a1���?̉��.v�@�{�z[	�f���2�K��{@����p��m9�	����\@o����Ԇ��'1���G��xu873�wfz���������2/l�e4��æ���\����@6[��	��Z�}޷�ˉ�PEH�j]��:�B��'�P�?��Л��B�>q���?�dƀ����!n�_��Mvޙ�QM�e���&�����B�ʭc9�o�a�=�DR�=��ĵ�P�*�w`"���Ɯ�VK�5vВ�|z"�F�r����)�ɦ�y9�8��l�/�d�¼�����}b[�v��&�@�|ڪ��≯�+>�iI���*�~U��(Q�����߈"I����z�mdE-�߷�9�+�s�4?��J�cj�C!�Z��@=���V^m���r�7W�8����[[�B��䃇\���� 8��!��ڶ�Ղ3=}��� ���N[Nٝ�Eʼo`�K���ٞ�i���/fK�X�ц�Fr�	���Ӏ��<nhg�H��1������	[:nx���Y8�V|���c6��g.�|+E��1HѹC#Bc���M9B�~�� ��"3:�tWuV��V�ҋ7����i�QD�M�Q��������a�R�Q#�A��7�rtZ��;2�^�靬?�P3@�N��	�&/������Z٤�Y}0���r�b�l�,�?�^�}��3�w�B��ާ�\�b��׃~<�l%B' ��(�-�����nf��a��y��_�]q/���H4î�:��1��)t0=*V����MݷKs̊=4�>�*+���M]�6�X.4BV���_{*���|z)�4�@��R*���i�����_�ݓ�����W��d�sw��ɧ��CF�F��`u�利*�s�iU�W"<�$�zm�"��M	x��YU��ۦ�+�{��4u���we⎅G�ޞ��[N�
T�q�r�>�w�),���z����"���%����_�����(�%�u�0;���F���~��(�4������� ��_o%aO2�����L�i�N?5���Qn�.V ���I�Ub����^�<����Y�������'�a`��2��/��Q��Ĝ��ۑ⺔>8]M5J��:��b�E�u���i��[�����ı? ��?#��K�&����'�Oy��.r3ԅ��	ze)���+�������q�gV�rvr��.�tx���J]s�a�*�
��\U��¦i|��,�K5��$��>!�h	A�r/13��p�R����'����hB��$j�
���uy��z��#�1�h�R��� �l�>��7���r��,<�<�mҒ}0��0���[b����}f��?���g���1����u"%#�H(M�dx�Ң1��J�a���0z+���@��1�6�L>3��t O�/҇y!u0-F�V%D.Ń��|��He֕.r
�Տ̩�1�qN�OR�Ĕu=�����hP�����3�J�Z��yb���D��לZ�sL3�@"�B�%z^�s��A�X$�q�C�U�l5Gz|�������p?cD���7T��� �Bt7�����{E>�l�V$�^��U�3O�d��=�C.r6%j��{r�Yg���o��j5F7ß��l�>�M+N,�I�Vt�>m�m���p�J]��; ?���$��d�_E��3�i>Fv�T��xq̩%��H�Wz�e\���D+�H�O�n	Iu�8���*��K�1�W�i^�l��X�K����q�_e���� ���{�{�}��|�6Q�������#02pMs#����5�bo��k��f$9��UXpT��7�x��d8+S����-F��C8�5nh�0�@��T�9)�q^����A�?��.c�hX����ߜ$Z�>|ֈZe 5[�Ǿ��G	T�;�uҋ�wD��)"}������SHT|�M�z:�;�F��H�u,���w�3�x����a���B/�����7"#�}�ƹ�������P�ؔ��\=��:f
�b�RK�)�-4|g��H���ʑ-?h&-�s�1 v��������W޵R{��Cj^�BE/�M�2A�/�ߐ��<ņ1��ǐ�-Q���@�g�w�~��ˤ��N�Su"�2�d¢S�k�G[&��U��M��I��������5}w��{G΁KV����5�Uc�t��U�B�9�t��L @��@��B/!������^�)��a|��8�?}^6�.�D���fĿ����ƥ�,~; ��6�}j��&��b�z'^��*���U�j�K?�;�&ӏ�["\n���G��X>iS��������n+h�j����f�s@&��kQdm�q��VD��й�h�Z��sPʙ�q�|)&ō��qe���ehCr�xg�&��I/拞��n��|n���:ǰ�YP�^HK�F�����V�hr~]Cބ'���ј�;�dABer��+%8'=�\��8�;/�s�V��ֳ�ZC�pD�W{�ߖ�S*L����Ȝ�I�U���~E�����`
�N�E
4�Tg4I��܅�u��mm�x^G�Ҹ�;�㔵�P ~�e��-&gs���0��� V��q8ؾ�߇|y��T�����nU�(ݱc]��I�<����$ ��A�xdM��C�%f��s�N0m<�:�1�TM|�<a�8SЎ	7�;t��4��=tV>q����@3й,'ȶu��[_7��H����]���c���b�-�5rt3tc����B���(aR20����ش3�ɻO��Kmm� Ə���lK=�kƻ��W��㒈z���$�;a�F��C�G�CRB-K�^?'60#�w ���R�U���A�.*uz��K����\4+�rE��qb�=�����c�5�n#+s&&�X��C�a���<�DL�!����Mt
��c�v}��X�&�ݨ2��2���g��)��P���t��6�����h1>�F�w:❇i�X���a<C*��w�9B���cQ�;d*A��w��L�_�(�[$7����X��=;,Z��#�1�jv�J�igr���!�'��fO�MZB�e'���A��E�k����Gy��pmdb�JGsj�Th���:�د��?�<�&|S1�LQ^�Q\_��T��u��gҎ��#�݌��-�A�X��������3��* v�̧���V$R������s��0��`�j'��3j�R�0v��b��ږ���_���ZDZtm5D��C!�<O��d~w{�]"�T�07�ni�'����Y�b�&[Y���"�0t��>�!�;�y�M��$j7?��t��o=M��T^��,��dM#�6a��7� Ix�/��C����Ա��D	JTQ���
�Bhr��XtQ�w"O`����xK��2¢(��� C8�؏��ד��G"�����ǐ���P��j-�4�_��^I�?ag�L3���F�6�DiG��.3;c};�VCz��?F'p���g<U������}TĘ)��+9�3�t�Ωk�OY�fGdPbM�c��g>n��tkdx�k{��WT��\���o�(����Co�2GB���Ϋ�t��r4_�7�[��.����.�V��G��:�\� s$/���*�^A����Y<�qM�p��M�z�Īg�vy�z��kq��'T0ţe.�hoc�� �|�Q+��͓3y�@�`r�i�<��~��%�m8' �1��L(Ӡ������V���[ ��'P����v�>5I^��ޣ6� ��m<��#��
��į��M�Tc-쒜��Uw�G{��|﷚ğ��Ei���+A#f�`;̗T��64sK,������R�D�:/�j�K��:Z_l6����*و���}�����!<���;ڪ=���|�Ժ\P�<i9�v�å���Q�3Җ6��h���+�A���]�|�o���}��;lNZ2\��n�j���4p���t�C�5��8��S]�Ӕ�s���{��$���o���j_~|�zc2_���S��؏\C�w���e)H��M.y}��5���7�6B��Qts%�VWy{�9N�2|�Rd�N�z> ޖa��C��K�ⴛ�'����7⾶�e�]GL�պ	j/��m���ϢE�$��0q�Bݴ;h��:�KE�������tخ�U�'�?W��kYU2p3�vL:��EhI��n͞u)У�Rr�/���CCD�5>b������8�/�s/�S��!W77D��c��8s|��4uB�9���e+٪zw�\9k��~T�_�&q�b=l��L�hY�)f�5ڢ���i�vXϚ��a�SXx0ϖ{zI�M���,G9�o���o��<�������o ��Ed�+zҲDz7�Ծ���Ir���܁bs����0ɼ�M϶�ڐ�E�IP<�Η7�=h�[�.������� "���b#��Z�D�<���/�"8[{7�М{���S�s��<����?d�s�.���^��J�4��FKe�� R���0#��Eu�{]�Y���_�ڬ�p]	},�$���GO��#��m`���(���Ǥ�0Vp��ǤpP�Z � ��P�}��Db�~��(u?���{��	�$�2ۍ��d"�i��sm{�Hcڞ�@�=���g��Q����~�W�L�f9�(�`��`Q[� *q��������v5�e&�[v�T>�ޣ�O���I�}�b��}λ�=�  S&:�u���,@���_G��NX �:��ǴX)`����B�;aV�Ft�2��1R���������3�W(V�"'%G�H~At�=�u�ݫn�,�RnS�i��7�I�һ�Izo\��!��G�*�'n�������[����x��\�d{��r|F�"Lj�'���A3�?�V�ף
uk�F=��n;���3�8G��ܾ��}�T�q���)g��#�zKC}���
cx��K�W'�P�N�W�n��>��w��T�1`�*GV��Ol����,�-s�	��in\J���_h��M�@o�I�洸ңfw`v&��.�����Y�)���~�w�@b��W�p�%/��@{R=�˂�IB���������.���Fb����iQ5�����Vy폕����v}L�҄�U�d/���Kq����"�����c�v����Pm,���q�^3���nJ��Po��03��ApNqڈ:B3a����bv'C\��;sg�-㨲Ҁcc;H�t��MN}����{�%LF��e����h�d3��Cz�M��lU��V�x&���nۙ��y�!=����a�[N�۹�����J!�!�zZ����*�)Lv.*0�,	G��Ss�L"C������B�Y�xDބQ,�J�C�oO)\<��h����~��)�gk������)�q�D��b5~��W�cS�[��L�i���U^UęE�5����xpe��d��V�U�Gh�hĢ�xi�������Z����%���/]}Qǽ&���]3.�`E);S��W��c��`X���)z��Jy����&��[��c���uS��}��������:�tك"�@j��-"N=бy�_�Y#��m�ՙ�����L�a���z����A=5Uh�`�R\(K�v3ϼ��fͪ�2n	N������2h��+�.:pƓAq���|��Ӗ�Jt>�L'�e��H��eP=5����%Q�=u�fc|�����bg�(2�֧4��r���)��ʹ�!C�u��>x� �6�I�Ӥ��dnq*��DW_�y��TB�x�'�(Z�k��A̾� D!�A@#��%q����)��ŖQ���U�H3[E�A�Ր��hlU��ay�'�B���H�M��B!g�&G�6:�0��ߡ$G:��bd��`h��ys�kYٺyMUr�$���P@�`�x�q��,��cI����k����Nr�M�,�����I�^|����@&�5�;���c�@&�Es5�q�0x.��왔�@�³i.��_� ?�C��_�~_�&<� 9�a�G�TX�8�#��q����P���ՕD���S��n7�$y�~�<rkL����I�8{	m_Ȑ}�ߥ���lH�e����RL9M[c����TN��Q�O��2?J��|q�Pɦ��w�ljX}��-�:��>rL)��Lt_*<���X�Eߗ���2\�j�IK���6��SӴ��bؿ�)��ARY��_�����ϧ8�]I��~�M]�J��@B<�3K�?&קO���j�C���\rh��v�*0����i���[D�<�9�E#��K5��r��\�7����W�3Ў��Sz�Mo�$8�,��?�i��׎�ᚯ��)�h�C�pӀ������p��O��M���Z��Y�RΩZ�VRߝM�-nת�<,x�I�����b����<�%=�%*\~��ȉ8�)�^w<����U���S�5�|:^���Jz�O�Av�8����P��KD�F���}AQw'���Է�����l�@��Wj�<��%jNЉ�J�wJG���\_5"4.�/�D�6<���犡H&fO��Ě
�~�%�zy���HSDj�]9�eb7A�q^>m�RN*0�#B���X`�|�#������WrEK����n]Syo�t/� ��vt�M�gn^H�������Z��P�����Ϩ����Fb�ӱ ]Z����լ.=��O+k��Jsh����8
ez� k��d�~U�Ճ����֧:(1��JV�c��Tm�o��~��|?��Rg��ˊ��{9f��#PprL@'�݌�rG��Ve,� �zdx4
c�x�־���htum鄼έ�9v)ͥ��Ԩ��C0�vr(rK�m��?���S����;jJR���ش�H��yWs&��Fp��89����	�O�έ�^��p����E�Q>%v@o�V|&˗�܏~��e��X�"�*A�.kC=���Ƕ<粦G����5��b�����g!z�{�M�D�ܺz^�Q�^�a�!oU�ã��X��c�7{W�,�P��B�\B(�����o��g�S��»�4��Htc�9�jP�c'\�W�XF�w�v�[��GO���Y�T�
:jb�Z�ŚX/���������UQ5kѹo!~�����=����Ω#�"4d�����,7��5s�"Lܴ}&�g�L�>K��ːe�F����\i�+	�u7~�;�����Srf�B���u�8PNk���� \�%�*��	�	�-+������0H;b��I7klq��uF��v��Ua���B��84}?�J"P^���Le�t��"?��܎�4.�x�����S�th0����TC2x׉cF���tL���A��,���a�N�m����[�P)ѧ�q�|JD�E����D���k��]��~�#	uP�w04�@����I0���+��9,g^�����e���b@��� ���y6��Û�漵�y"� 4��;P���mE(,E�h����zxڡI*a�F�}6M���	/�6��7�OMmj,@�U�9?7�}����>Er��2�ȁ64�@jM��asG<G�R�Gz�\��� ���1J �r�?%J�T�"�̾��!ZR�;�vm}x�`]LK/�A��Bx1*��9��N�P�0�!�Xtb������G�H��9v,�pL��!�8
� �p�� T�˳��P�B5�$���3.<S��c�Z,).��#m�=�CB�d2��5�L"-f]��)���f�_��*k	I9j�@�X86j�<6c��C��N�{��T>��U	����&,j٘�q��u�8��_}
@�i`�U�P�?hC�pt+�k��	����S�� �gr��{�/e�AE�,���.״1����������q��m �0�Ov�eK�#��M����a�ǋ.�xJ{��y_6�v9� l�C��FE�r���M�'xX��K6a��:���%��LO;E���7�S��)������Z]X�2"��שm�ʍK�;�}E�SSVn������o�D͏�Y�a���Dv�U�ܖ�b��S^];�pã���59v`��%��!��+H� �h�2RE��s�>���B!v����m��a�'�HpwDqA�������"���k��l�?H��:�lP��/z��nZ�5\s�u��Z�#TA8���X�)�%�ڂ��z����8l�_�zڜ9YB7�ХJ0�|d��4��Ƹ��c���@��bk�G�T����k���j��֋PU��I�DJ0�H�FW��>�]����7/�t��|���t؂o1��[t��=-�^�F�X0�b�~�G��]IC.;��aһ��oq(o�,]��0'J��Z�dD�����h��y��ѯG��3n-�溺�a�F�5/�MYO����7�����Jw�3՞�ޫ5�������LW�;ï�������� Dl��\R]�����h�$�p�<	Z_s�[���_@�]`��P�]�j��Z�qӝuK��w�f�uŝ��`�1��N���-M%x[?�[��sq�E���o�,�	��N���Ñ[�S8���3e��_�ԥ����bHR�NV� �1��}�@
�`��fn��K�_'����EE�G�2�����N�ʖ�?GQ���Y���L�zjMv��T*]9E��N�K��)�%�� ��D�:4�(l������X�����0��4��YݺL.rm�_�����Q���i�f�?օ�@2�r��;&b-�� ���jxp-�qg����<]�J�U��&	3��#�>����ѨuA8��PX�k�o�cv���*�M�u�b���R!&�� �sa$fd[� ����:X�+�4:,���D�����C
�;��Oť�[dN��g��.̑䮢L��&k���U�7�����c�Pew��0�{�C��kn���]j����/:�2A%����' ����͐�[·��� ��U5��.��HZ�w��9Z3�ü��B�r��'�K6����f�o�1T]B}@��$ؑH���i
��T���N��E�;�R�^ڞj��?�`yk��r����ETB�&�P�s�B������\t޴�'�0�mϦ5큷J~�q'n�y4N#��G}�J���j�]�lZF��i5@�;=�f�i����)}2�-3�V�Ah�U�7�1 (�D��>�3aZf���x��� �.-�����#z�S�~��9#�uFD%���q\)�O��-�|Pׂ=j��D=	tF	}��-���k��뜞�^mE���ł�8�n���J{Ŕ;N\ף9�SR����r5^C'K�/֭�1�R5"� As�3T̱htɇ�� �=R���uV��6�ѝ��0|0��F5�1����V��{�2��j-�
���'�W�������U*�f.�8�Ԫь�TJmeÈz#u��2Pm�^��]��*ɇl![Cʵ;���+S�>Ó��+AZ�=�c^A��n�پ*�@�]%m�3շ��F=�1�>�� ����K��в垷��w�G�I3�,01P�ޒ�Ɓʩ�s�T�>�6��^.|�
)/�Hfs"��ō�-��H��:��6\< �]�rJ�15�EM��_�n(s��k�7�[jHmOζ��(�;�M��`�	��M^2t=l1�Qr�Ûh(]��WɁ5�����b%���<�؃j��5���<{���n�/�*=(����V�9�b�,�ǎ���ax@YV��������%k7��8%ψ�Y���6��į�pV����ߣ% �7���Z��'BS(��X�)��]i��s����9���_�5��<W����ziV��son��2�7	Q>҈����B����CG����y�b��w�S���	a�s�e�~��v"�߸~�n`���˗__��s`}h���U�==�ޮN��z";��q�e��Um�ȫE{�PE�6V��+v
�L���WFL�e�;`S�M/ZХJGs ���{�.�u�xQq].C�w�8�M�R�o�~�Td�k &[���Q��B���Ϥ�������jߗݷ�dІs���<{�W9$���6T�v��I�'U.������j֞�������F#Y�Ct�1E2�f��A#�6L��Z\=?��j����v�N~J;}7�L ��)J��m4]���sT��f�;?���^)I�]��ʡ�'6�4�d��`��Gk�Zv�	�@L��bpYIyF����!�4��2���f�h�{wэP�Z�	�-�#��_�;ZHm���%;h�)Q��|؊�3��&�a�I;��8tGxA����mj� x��K�s$��f���xW�/t������.$r�INZ���p�0��S�B)	�eD�s˘!��N��Lr��P����v�3�7���h>��(�H?ɖ����ȹ�~zE�>���R^���Jol�1Z&[2@(FZ>����d6֫s� C}#P�`'}������ӂ�:���0�_�4Py���m�:��ā�lK��'���:�dUO�@���U��W��[q�Y�i@�ׇ&~�ɝb\WQ�65ߚRLm�� �$��΁��n��u�L��%?S	VC�����-r�5���6�Eo�;��Y�3PĲ�J�S�+�ܧa o��������Ĥbn	i{�mT#��!��3x(���&�X�2���9����1�[>�M����"�p�MP�9px���Y,����L2ك���	Un?�_M������H���H�Ut%x
~�}���\l8��P��'L<��h�&��'˗�>�Ē�԰��8'Z]G@ɱ��v�����@h(�y��ԅ&�&㉌�i��B
ً[��o�@����M>��s��BZ:v"�����Rtr�.�sjK��(�dvV1�[�-"z�h���ߘc'�4���[��~	�l�iu�gR�*����F��"���	����".t}��%��+��yb�����nd��ⴧ���;^�e�m�� �'��&)�u��/J���oGE�#8�� V�c9�C�S���=Z�O!��S�����K�!�M�E�|��4�lo�욁�y���h1���K�HNK;�'<n��;��sN4ĺ����25խ�/-j_W��2^��ûb5�M�vܑ}мV��X���U�&8z��5�֩�PRh���F���^�s�����������o�@�*0�U�'}M3ĵ���^{�ZFt(:���s{����2o�	��e|�i����o��lҧ�xY2q2v?��g��҉x �Z^D�&����\��t���|y�?E��6#^�J���hbH@���V��K�L����D�·�*@����K������6��T0�aR�3X������~v��͈;R ��V�5*�ݞX�)*$f�`�����m�k[�E߾(���G|�S�0^��H�xTO�5��3�^�Ծ8��U�6{��4iQL�<�jAn�%O|�4N!���%�NԟrC�C��ť������܇&voɰ�����by�`D	I^TeHLy#R@��<2(�ج��8�Ft\�/+9���G�=3$�N%��5�CG$�����P�O��cs�Xܑ�؝O�����PR�}'�*;;O�$���{Q��n����@���f�]w�σ�l�7�aFy�2�����1�)��e��>�;�9�R	��z�rG��ҳ�/���t���)`�ky%�����Ch�!m�����b������Nw�N�G�3�6���q��ޮ��`BP�Q���~ʻ�-��,��)��71@'&�uS	U��&n�f ^>����P����3m;�)b�J�^i�Q-�[I���+�t�v�^Hr12M���������o�)��7S����a�X�$ƅ:���@���oG ��_� }�ԁ��g0 ��3�x�r���Q2u��H�ݻ�u�?C�Y�̅�~�#X�.��?�+g�Ex��E �6�wnSE��9�j� � -�*����Q�U��kiI�Al`}2��R\��-�p��e�n{	�*�(����f���t>D�ct�M*L8ԑvH�7�$W�^�'58[{��D���,��"W,q���'J�g���q4�.�	T����j2������	�F'�����_"����{V<�4�M&1��rN������)K��Ѷxu�����+�wB׾����Қ`<�Z��e�Wх� �@�Z�}�ҷG/y]|�G��
��C�������(�[�u��p`�.���;!4n�ᶽ����ϖ(9L� ����-(��M/��py�;a����(�e,W�X�b��ֳ�p��[N]����Xn
�סR�u�bZ��o~^@�>;q�b5�:�A]<\�6�U����lȲ�l^����[���ّ�%��AB�Nϣ�����(�n�<�>�BKa�?��a8�T��>Ip�v���ԏ�e�#��R�h4��Xx�(�4�x�8�iϚ׃��^������7N�����-��-&M��W4U�L6���D�Q��P�j�E�����?�V۫K�S�Ӽ���u�{�WD�����|]���y���s 4�E0�[��4,.sGI���>1y[ç��?j�rVnmݹ�A�B��k0HRcC�*zi��T�&��#�u�!��D���J�0V�w�� �G�u/$<�#���ff:"�RQ�>����ף��?��3�^<��c�dkx ;*7qto��e�a��W���g>�\�P��G\e��9�Ę$����֕n�7(����>�(h�Q�V��5B\(	(3�=Ɛ�SN�!((�UXM���o���C:��AZ�]8�K}`GdY�r\~���?�a{ѝ�������v���� 8TJ��i�1y-a��M��,��9��=� <�	���I�:�j)�ܢV�_f�^�ӸOo���X�bh�-Q@�����@��[��q�'�A�\Y�8��D��Cݪ��4�qG���ڸ�:!����-5��T-o뇭��r�1�%��܂��ii{���f�̯��BX�1��*k�ЖX�8�I0� ��Ĵvb(*�.�<�_��7���%Km�����e�wQ*��nJk���J��p0�]�X+�~2˨�x��\R�C��Y���ݤ8۠��yϡ��kLN�t�|N��4	H"j\�V���3ޮ�˱Z���Ӷ.�Z�V�`������..���Uf�1`Y���Q"��v��^P�=�[+ݒw��\�?�3塂����RXf`�cx�<\4��H>q���'c�������ͩ`(S	�ᥰ1��Y�#��OwS"�S�e��R�A5���B��OQdL�%iW#�ֵ�$:$�N�׭}�c��|n��^WCH���m#tÈp�E)D�:6b�0���}/�Y^�O|��(w�]�K�ΠЄ�@�lM)-.Jx��^��<�vEǿW�#~q����he>A�@m�B֞.�n}D�E,0Z���H��|��>T�N%g]4�!��Z�C���@�:ۺY���_澦gPa-Bw%�~�ꀸ!�qA�B:�qC�d�� �e���~�����A�I�[��P�+?Vk�a?(�º�3��{�8oШ;o0��f��cw�K�)z��@�jen��Н�?V�f�l��P�|�}P�'�[��<���tj�&����OZ4�>�ܐ1�����j�J�����ޗ,RC��6����H�u�P��],8�j��<��X< I�u�L6D���d�t�d[�il��O`��08I��ظT��Ve"J��h^1�j�X�p�SC)�o�=.O��$�+��X�&�顢$
�Sꁁߟc]%m�x#pD���®�,񌎰J�a�a��Bl%��0̖>�%Ý��1,$1Д�X�_�$\dO�-����PҸ�Y�`UT7s��-)�rg#vvg��c7ⲥr�"N{��V�L��tAvOq�0����<BH�Ԝ�zy�*=�BN����X�_J߬���"������cѢ�EW�[��3�����R�?�����1L�d�C����1�Ȅp�(#č7;_|Pk*��Y9
���'Pa��N�Z$Տ�yս �P�x_��|� �L�
���$�7y����p��a��v+����iv�wp*<� ��,U�e��e�vγ�1�W &���2�2��t]F��)/���b�~r"�!R��.��NB��ȭ*�-��`���I
�!1ܣĩ�J��*��Ϩ�k� ���6�{_��Zg��gW02�RQ�D�[�����hFX~ƴ����.��p;C\���z��Q�2^���>[W�S+��L~�y�i�k\ήj����k-�]��R������bs���zD����剋��C�u�y&I�"�j򟽸����U	��!i����1�]�7�����?u�S{���nE 3�rP����'��(���z�\��g�.,���$ ����pP8&�k`=f��/�}��87�2��(o�F�>L`̒�ndr�FuSy�Q���	d+ �ȹȎ��^��O�xdU^S0�?�����ۏux��FW^ ͗���b��m�ZU��"��gT�O�p�~�Jx���9�I3����8���:!2�<\�v�z�$\�i71
Ibsxh�ݢv3~Fֹ�� ���.�R�����u�$�;�02ܗ�Q�0.����8P��z���0�4$�4���:�׷�n� H7��K^�$Ӂ���O�Xݘv��d�sݘ��ٶ���9��F�Gq�uܹ���\�@��|�͖j.NL!�<�(",����(��Fň$Vǘ-�wǉ0�����1�f��5��h;6&�P�Xe�X�s��,�Ͻj
���f4W�ڊ���K�
�qx���MɚkܷM�"rm��m������,a��Q�8ypj�k�D���aU`ɥ�&�!IU������e�'�4�6Y��Ek���|}C�`S����a���n;g���p�,w���8���JN�>bs����n�I)M�Tė���k�
��6a��=P.�!��ng���?�bR[Ʀ5$�G���k�,l[�*���.D�]�ftV�&��}K��������,Q��Z��PW�9�3+�nTϮ���~9h��'N\.3����ۚ���d��f����e\�ߑ2��W��r�g�>�L.�ql���>��A������w���<,�˱g����m���i�e�j�1��S��2��p2��xI4w�њ��\���}\�sr`�	�6�:{�&� �,�^3��B��]|Q�@�a�D
�%?5��q�U���KY�����7��[�'	1��3�����rU������DjOփ�Y��aA?�He#�{����f&��c��Y;��y�N�|U�}6Z�/�[�=ѓfð��#c�5t�������{$� �Ǔe���Y>���r�SKv`��No��UӝD�x�T�}�3С[*ڐD��'i��MI�V�0Ҫ����`��F���Zd�tk�fAg�Q]X�!L.�2:��d�m\��nA�KH�oy��|�Ff�-4"�=	J�m#7���7�
ݿ���xh0ɴ	��q9<�j������!5�����-�pޛ6j����'�]�ׯd:Z+�����.��f�(*��ś�������O8��l�%q���o���Ϥ2�WI��4n�'��1O�Z�T<��ࣂ����e���'�g�3 �p�^�אSV��<�ŝ��'���Y@9']uF��Hݬ�� �:N`DL��jc����
�b�bf�f�wm�u"S�ϓ��@ҔN���d	��a�w��^��J��7����0S�)�ީ�����_�;�kJzk�x#u΄�hzG.��wlo��3O�o�'5q�`sn�n����k�Z�B��&H�PSCXN6rO�f{#a���r%�V�ȫE����&is&�G����	�X6�Y�b<P�Zfg�j��-�@oȑܺ��P�6]��oK-����k<���Ӊ,S���}�\���zz��څ�E��M�\r�`��wq��C;bRӢ�X�ux &��-%H��~S�C ��2@G��S҇��A9-�}\'��0���%����4y$�1b����Ce����F�ã-�T�3��Vg�Rk�w=���k��R@R�,�����u5y��H��U·�R��#�����uau$n~�M$��mj!�3����|�z�|�u�ϹH9-*�S�D�  ���]i��?��V��]�O��\�]s��ͣ���d$�����{��dn\�8}#M[���,�#����F���_H�:	J釨��6��"�̘8�ۼ�|bG��1*�>����OԨ�|%�Cڙ
��(�zWg��RVi
��Xȫ�>&�� �VRz��,q��mR<Hɵ9M�d3G��g�]�y��0XɃ�>�m�Rk#��,�o�*n�	�60C�׵�m̹�7�2���Wp�
#�L�W���j�NO
%u�&W��,Ϗ�sk��7쒓���.85r0��$3�7KP����J�`ĹI�����-��36��ȵ6J��Ѕg= �"��B�_'�n�«���#U:U�7���
 d?�?����#�����Gө�m#�d���|E�Ra�%	�iY��i�a��k;�j��p-6�6���b����'sSm�[����#p�e�I�6q���m"�[*�&����6��ḗ��z��NUħ��>����Uh����4ݫ
�;l�\ 5�p������2�O�(�R�f�8w��w����Sj�Qr<��h4���	�ۻ�A�V�3/�f�h�*G��}���-��O�����2��Јk���T�&v�68������}��`���2l5z�s0��4��m����',�''2DأŮ�^5��bΛlΎ�x!Lie�ɩ�t�{^�ňB��v��rĳ��ya���VN�3u5��ϸ4�]#=T�C^�[��>p;�k��G"�?~/f
��h[��}%X��c�R�u����q�ܦ?�����LS�}EFqr;ʜ_D��ڷ������^�].:�xX_��fh��U*���Nӏ�R#<W���ϜGJ|�6r�q@]@:A`����z��E��v9�����1:��%�%�B�{bC6�;E���M8��j"��V*P�c�{��x���X8y�?�o���PJn����n=�`�����;�������:J�����B��Tu���iF�p��˫9C�����|_i"�wn�7ޜ�.US��KGCP}fy"Ţ��w����$lc�
��MyC�~&���@w�3%"(�=����~G͸��������AB�dЙQ-����� C�:Nh���xg�K�=`�P^>,�����X��"��k��[���w��?X
N�La�r?���<m)���^���W�`�DOt����(#��kyr��d���9\�
����ʔ����G��Gl𑌊_�!�=A�:�����߷�U�Ǜ���SY a�6�ؗ2�]�����c?����~�]�ƛ/�M�?hCQ?N��Y"t؟	C�,{,�&�D<�ߨk��x	���G�1`�X����ȽL����9�Cc���1
�o�=ql�Y�[�ya|V�l�"����WV9'���vp��3b-�@rH���	�̻���A��������>��v�]��V�>�?vh�+��se(n嬿�)x���9�2*�,,��-Y�Y�D�4Sm6Uڠ䓣��D3x�}�,�4*oI�}$��G<��g�*�]V
0�tA�>��mk�&��Q���5�ڷ���8��w��B��i�Dᘒ�l�M��� #IQ�H��&�C`�VF�we[~���4������^��z�Rn�A�*�#�2�����>�0#Z�+�̵��0U��`�mo�R�6���۬�ѵ�[�Ŀ��݅�e:�2~�t����ٹ�Ѕ�`+eB	}�Ϯ�_7���@������BѢ\��袖�% ��ެ���Y'?�M�!��_��&�T(�ΊJN�(�����8`�k����gFG���~�J�A����;���
y ��ge�O@��]Z�����os�P`Ng��sEa�0�O�GZ}���^����=vK�"W����x�?m��ơb8���bR漗����5a]N=���E��q�&� ���L��e���XCkq���$��tV���Z0G��Gi��	�K�\��%3�9W����Uņ.$�
������/1�.n��^	�3�W��>	�C�c�\D�p��7��ą1'?e]�-��ʇ>�P�\O1�Yp��^� �|�����s,�ڋ�r��ϛy�*�9
���a/V��ە�W���X]�(V37N�9�U��m�4�3$�'����`r�4
���Q�=���'�x-m�DYdS�s����o����L�oŽR^�hH8�6qHc�̔C.j�OX��I��p�ڳc�*��S�	�������'&�b0 �HD�v�Ϻ)�8��+�l}��Lm��r�<ԡ�䥹㌕�	��r��{�+��wlI���:	B�P�t�Ua�8�znpQTn�!��5~E�P&����v]�4����z��\����\���v,�[�<�~Y)���?������\+�z驔�Җ���RYů�̗C��e� p�����Kۗugt������l���όS�oNuc	�����#�6�4g�'�zLV 7�O��#���"�♛�zG����=Q�5���@GMm� ,U0>ſ��0O�c#�I8��G2nG�s�Įk�tH}R�ߎ-ϳn�]!Ď�q�f	��H�Qu)0��$%��H-M]"�]B��!�-�Yz&��X��#���_d� 5���IT�������8wE�y��k�7_�����&X���4�>�>����������Ȋ��a�'�菚&���s�?���힥E�7�D�[4��<��КR/e�f�#����\���u���i痢�6)^�+��p�>��me�`I����gEd���x�gKV͎'��N���W�����zx"qLf�v��SF<�	������d �Ǆh�ʨw ���v�0��S���J�0Yf"V$=[j軪k�v��hvβ�(1/��M3�f�	�BO�J�T�׫�l��+!%�F�p�/H|0�l��\[�Ho��b'K@�G���:��'��A/�l$9�ɝ��87I̪G��{��g��8}�r����|��R�Ӝ/�J��00d$Px]U�e�?����!u�m���ܳz�G �)L��xʉ�%�<t�$��T�䄊g{��8j����|�.،Cd�f�h��wt`(�.���W������t�%��J�h�1$[zK�ϡ��J�[�X��' p�۔_��gas�r�`I)��ծ�`}&����L�@��ݗ��d�r���DI����l����Q뜟xf�F�<��L);��-���j??�B����R�=Z5�+���������%QE�Us����J3O�\�I�N�H�А�"�}�R�aMk�'���%�c����~�1� ��6Q	\�Es�/���[؅����\�l���6�l�V��	�<U���fpA?NI��d �	��U��L�j��'>"���Y�����&s`�������ޥą
�@�ab�xt�߿?&�<����A%t�u�ju�g�b3Tj2�����X��`ۮ�t�*:�Uat���&�V";*�%��_�jd�_�ψ�JP����X@�SF��!r�H�eC)�	t�r|���^�����l�A�r`
��J+Q��٨�T�,XU�����<�tl��i���x�߷'Q1U��A�t��K#��o��oU-M&͝D[_[�e8?Ֆ5��;�_�8�Z$�b�?��0�O�P��^&�=f�g�s������pۇ�f��T�O�,&v�f}C[dsl�T��l;
�����Kr�4��lϨE����[}	?E-D�Y�v���@]�%Q���#p�j���2!�M�rQ��*5J����r��w,q��g7[��k�*,Z����k"1H�p�YE7* *3�ܛ�6�g/���<[���:3`W���BQ��o�^S�Z}��S���9�rr�����\��g��`��L��VF�f� ɚ��SmE%�yO�e7��/y�r�����6{s����M��
8�%R��Y��%��"�b·,�G��ÍYU(bOr<6�ǬO����m!�����NPL��yM��b;���7�e��L~�Yk�]�M 2� ��̵_m$����m�࿃z]N۶���w%#��*�"p8YsAAb���C��rq�P+���a.r���)��$�Ժȅ�I��Q���~a�l�n/�����[�a��Ӥ���}12�QT�٪p-����YB� �q��&-Tk��e%�
C2�i�V�EW�xN�>C����u��.qRbO M�	Ɖx9��Y�!�P�ALw��{�\T��ޏ@L�v�#�>���2~�2.g�һ�Z����9�p��	�_Y�<t9��'� o�U7"$���w��ΗM��3���H��GT��(�G�~4����1�=���.�ؽS�!d6���0��5��@�[<�,#��,����
�����v�( ,�hX7U��Z�Cz$8�~��2�s�˨��>΂Q�{�ɒc}�ҹ�&��������,+G�|+��=�S2�C'��p�~ј��0�p=�����q��'�[�(�E��q�>4OY��ُ�:�8�bU�DV�J��яG��f$�%���g����t�Aٙ�)��&�+^�\c���	"�N�p3�c���l�쐷�&��b�#�_ =[z^s �f�%F�:����x�C���Ҟt_�s�5+��Mg5��N�g��P_�i4\I#^M�.�qSh��o��	��"�%B�@%��#�Ȩ ��e��o���J��cԞ96�>�ü�7}�P�g�o�
�@׺���{�aDԾ'm�� a*���n5��]Ȋ�$}MLӄ}�~h;Jfu�Si�E����P�v>�M�p#I&8�$2�������ۥ�(A=a�:��I�MBs��S���^�<x�38��nM�ǹ)�ױ�x^
��V�P���������G�%+E�N���n�ȆD���F��D��D̻ ���m[!ev�W��3B8Z�=(�]2��]IvKpp0ހrI��`����7'�K�6*q�7�p�mPm�8�]_x�5���E	�!�ަ2�:a�ܸjPߙ�/@�{�0����U?©�)଀��RǬ��뢛P03�����TrQ%��w��B+����n& G��z��1�9���6B���2�3�v�)�h� �����Q0��
wټ�(W��� ��k�����M l$kҥ�h�� U��������g��U��,�N4�W��M�@�=x&n �����|�t���6�r&n� o�����d��s¿1��N� ���M�k�Q'�V�4��`-��L2��J�л�	��b��<|�SY��10��6�t`�)�2�ڽ��/�^dAX��B�y�����Ӗ��1�wu 
����ƥMO���v��<bs�1�RTskz�j(W��c����A@�@K�}e�c�G1�`��V��LW�U!�[V�g�ݰ}
�d�.��1c�*��|��<}�R�w�$E�^V��A7���*�����f�����CB�p��j�R�����kY��������m+�W|����|��-m%�C�I�I���4/��|� ��-�]�����h�s����鑩���u����n�_I'ҕ^��3ɑ�(��#��?ح��:a��j���R�rnL(Z\y�*Y'��e�4���s���V�y4j��(0�:Ν��!*|íq��������(Uuzist�%�չ�>_�Tзd��P���W�@�v�/Sr�H��x����f�b6���Q������ʉ��٫+�B'-��p�aߝOTΉ�EOh;�{�CG��/6 7E4�M� �/�l��:���j}�T����"��]��/�V����jp	��Z/��$��;"F��٪)��)����	2]_ǌ'��Z �����Z�_������u�_[�|
@E�S�zQ3o��IG�b���4k�ib�x�RK�[o/y�ƊIŪ}���%u;bj��YN�n\�9�#44��aː6�C�(�R:P�Y5+�e/�a�$��rT�͛�~U��!�?���A��"wK����R�G��x�4?�����������*���Icuδ���SJ�MiQ�#Y�$8 ������ٚۉ�ԥ?2��h�d�!x�� �WW�/��?v�F����pf-<21�E�dˤ&��yj��ݟ�;��)t��}Ifl9�1垓�9���i�!Ep%��6���.�I%,�Y�$l�0ͷB�d����|��G�P�ۼ녕�zz߄8���uL1��x(�v��5��*�/�ǧWrM)�5�����l(�m&Q��.��M��tbE������[��m�C��=�nA8�����b�����?;����&�($XԻ�5�>�	5�7A�ǈg��[�l)���M�?b}�+>-z����4�D��&����a��ʜ'Oټ�w�RPL|�~)��h����e[K�q��	X���پw��k�Q���nE�'zf$j].⁉H�m�Y�e	�]B�Y�Q�U�AX�j��p���ƣ�����Z���m��owMc�2Z�%a�{.ǐ��HrX���=Ib���r���ǝ�P����i���	Ij�|�� �S�鸱����&6�8|����f��|ݖ�ԁUZ�t�"���� O�G�Lxi��]��)aI�r�(�&BAD�Wg=Wr���F��8dv�����]kʔ�f�c��y�e[�PT�#U�OTO$�,�[r�5+������B�Y�K2Hs�㷖 }@���a3r�ggA��(���4B���ph�%����s��W��e ����z����4��1�ۈ��+�( O��nh'�>ŏ��r>R��-�Z<2HV�nƠ�a�	�L�UK��i��3���r����F�6e���$�y����!��5�3Ơ�a�K� 6��N�7F�2<��`�5>��<[Fs���=���a�}1dݷ8���8�(3(Ku�ػ��;����\�S�oXe���V�`�7Oh�4m��3�0��k�K��s*��htF?��$(c�V��z;ʱ'DQPF"�໋K7sS+I�MnwOL=�q$��{.Xf.��آ�a��F�f��^4�7�L��E�4� �'�3~c�;�NE|����d@u���פ��7�ρ�N1���~���"�����F���G^ӺתySc��q�`&����(���ۄִ%�̖�?(	@��$v�u��LP�d���d���ѫ.���>�?��X� ������ތ�R�	X0)bHC.ڧ���IR�M�32��(E�:vÕ$F2�G���bItЮɳ�f>���rNڃ�j�_DD���V��y�RDg��4�w/�+�RʠD���Sj<s'1�u)"���)1H�
%'3���ld��=�/��X�1TǬ���Q�eu��0QI��S!aw��h��!�Rxۯ~C�\F�8��qP�����[�V�����k�6� R�_�O$5�+�\Ԣ�V����DH�{4����4!��^V��l4R�}��
=�:�����n{�n�#��1�����rqí���>���-HdY$�2��K�v͏���"m;殎M����zP5a��J�b���;
�����:��Xb��g@�);����S��nS�H�Î�6��t(�8ʠ��
�����9�e�f���8ڜ��fm���,�Lq��I �1vN�h�R5gS�Y+?�4nr�Y�!{��-�����0�P"�5B��0~��Rs���A�:~�e���S�&�w��!#�ˠ+�½��R_7���q�yJj�)�����5b�xDA)ƴ��N���BN�#����GG8�K����ꉖR����G!��B�"��(�:����K��l�FR�ws�ga�����D6�@�
oݗt���������*�s��ị��f%^?���X�"[-ه	��{����%��e6�s�k��d�ϸڍ����2�!^A�f�X���4���Q���_�"^	F�TW]�V��}��?D���I���s�[F�[��]��QZcPl�hƢ�zh�8�R���&�jsP�?�T��e���!1����/�$p��@�]T��
Z>��?[���/~+�&z�`�$�|����Z�YA0����E����1��	e�L��ER�����p�'`��~�u��L J�,՟������#�����j�;�@\W?�в2��`J__�G3��2�=AJ5i�:x��=i�TTga�=ɫXA��I���:]r:Vfu �\� s{DT]@��`P�/:��i2&cr�(�Y�d�t�#,%&���W�>��(�g��#������/E�F+��V�["����A�P��0F!��S�0��A�6&��̳K����`([�N�� ����G�{���������%e}�����`�F�6N Fo+�����e���o��w���mmפֿe�
f8C��k�ů�6�[�,X؉ۣ�l���
��d1���l����|����^pj�I���]�e���=v�@��I}�X�!t�� ��Z$�_
�@K��j](�<�yǮ��G�T�]8��#����|l'F���w|�Ė��h"�1��X�X��us0"U��l���z�x�k����,�%�֣*��OīB���5�DV����ڎ���X��/�&�f�_��T�O-���&֒���t>gkw\���޴�]�h��(F����ⅳb!o�Ӆ�:��V���$��D������k�J�zQ�ox�޻C!��_"���Ɛ�+���R���h$C�9�c��S�-:1ni�ġ�)�Xj��%���(c*I�TK�z�s]��# ŧr9Z�
��Ke��PE��AW�}�������*J��z�j�0�K�.��~��`kVpCw��M��!d��B����Q�>)E��#��#R�XЌk0�4ݡ}�]~}Z��=�,1��c�$���V��G���I�4ϩ�y�L5��$����H��D}�WQI��R��m����Q�ƾc�OqU�s�K\~���~�}����(����ӏ�Q|=�T���c�=����P����eW���ݪV̡�@MIv��1T<?�~'GK`�;�tPI6΀��~���ȡ����U�n�e9���Fe��@0%�p��7�zl�x�e69k�<ˡ��1x��c%�|��>���6��"ǫ|��bdݫ�L���bH���N3���T���@�s#�F�K�)R&�d��07 ��<=&���q���;�C^��Ӊ˜���x�3-'ZYqlXR�h��������/dՙ�X�8�_fb�v�c�w�2�
�����9qntZ����^�|H���]�1> ��E��������;�p�:��f��X�=�&�H	j��`I�ۊ�W��UD;>�o��-�NF��c:�`��ܳ����}�6��E{�W�?1��q�"92n	i��8�Ԉ�������hd�ڃ	�	��QIۄȭ��T��6n��8��I/�?"'_,�����F�or���\WwZSO�%�A��xyE�:)JF��5���2V����D>���ѿ����n�]��A�ݕ��A�;K�z�)`�P-}!�2�-�P|8�B��l�C��I����K{|G|1��P�<�t����b��U)�m�N'p!�499t�ݠ�W�}I��d���N�쿧�4�Y���#������q��KFj����m���[,	1�ɪ�=�A-�pg��"�}Mc��⽊O�̶�>�ix��$YeL}6;j>i�ۦ�8�{r*��yv�@�1
 (+Y���i�"�*�7��ʜ�8_��E(< �8�6 �|�όH�5��ߛ����l��9zL��-lf�z����|�|,&˺z^�9��+(D�Ԥf�r#�{2wY���� ;�'�m�a�'�独�:nG�[�����������J-m�-��\jt�]l����R^,��N�i>�Ft�۸x��	 g4xV����4���_���='\X��9����3-�����Ӌ����Y���ϳ�����_�\ʙEw_�"�<-��Q�1�<�B�j�V�����`�&�j��A�����0����
ˉ�/�%�'p)s�s�
����kc홤�� �T�a���&�A��6(8uċ�M���?F�kBf�$y� �ˀ�'I�!�R�`)���J����g��Yxqo3���s�E^L�̄V��BA�����3؂z��Ǿ"�4��y)s̎q�^1�w�W�Sd���Nv���L!l,h
�g ��<�D_�7+]�k�hsj�{v}X��,k:D'
�J���Mg�����)�0���ɣ�F��N�V�B5&��h[�zD.AG����5� 4=D��������|C�Z�buh9��F9#Է4�� �?	i�;��kh����	*����f��^p�T�����S�-��l�=�Su��麌p��
cڣ���6��}"�#׺�<�Ց����$�7�����܌ynޠ08e�B������e�o�ho៴"���V>S���HR�PK����N�4���[�Bb�jsJ�e\�����!~���*NmI��R����ʻB����<�a�`��d��g%K�k���(��gaJ��%�����3�Df�'e��p��]����� 4�@��F4�s��"�})��HYs'���&m	(FD���R%ףe��� -�E�-�9u���:m|�tt"�lT�����/����� D���H�Q��P���P0��h�v�NT0|W�z�D�(E_�wƶ?������!į:	O����s܈j|M�(�`�֋���� �ƞoǅ��.B��e�0^���4�\�n�u���V2Lܮ�/���t�4B>�[��TdP���C�?i8�VV�n�"@��fGuN���՜^�l���"�����^��!���";��2m^��<�
r��V"�9�UL�J�q��y����5���h��S��"q���9K<��aDw�EY�Y��XD����9�*����:Kz+��y��L�_��&U��r$�� %���?��.��Y�4(�P|��*�����S�3PS�Fc\"�d�����{Ḽ���*�|щfW8O�덟�m��~׫T~n�)w���@��������^~`�X4�Ў439�0��m8��,���-`���+�H�r �K�r�5��Ϳ8|��,������ȿ�uA�:���ê���F��NV�Hf�H���C��A8�ƀ��9�0R[]���i(z�9�Qc$��	���g.�uTĎ��t�KU F��\�HQI!U��G�T�<�N��f�*`SD����QU��Y��K���OK$uq/mߟ��u���q8R��i����ܥ���j+��a�J�&�}�!�)Q����NlW�a�9�{�>�U��Ĩ6T�r����*T���EX�%L����Fc��-����9fSH�b�@��x�9|z�a���Θ����@�~�h�w� ���f����>ٻh����B�_�a_#�V[#���q�\�8�����
�G�x����j�ƒ����%��i�h��� Apv���)�'�
}|�m��1]vT
%����pM�H_h��z��D�� d�C�W�ʇ�ǽ�]�=��@w���wD��X���Z���%����A��M�pa�a>�|�[z��Ʈ��ڸ��f:��'ݷ���f=��_��fkX���h�!/!��ʩ��Vm�%�K�`����P�-���w�@�^id%N�os51�Q�nr�nd��M��:�e��,ˎc��L��������J�0��S��Br��KG����	 �(k�+<���e#Y�Ą1��~F��zǂ�UfBX��WJIc���D���_!%(�WK�}��p�D��9�!�����Pl��6'{rb&j��k����M^C�Ve���i�'���w��b��n������~	}�,=�8�I����݆2���Ν��^��靉� ��T�sL��V/f�ވV� eE0`,E�G���U����?�1�v��)�����!�3�t�������5�[Og-%�����H)�z|К�J(	x۩ר��h��[��˸�1 &i)�L9%i,���J�gR2���sw�n�f3����k��C��>([%H�y~ �y����촶0CyVI1.����X��I����^)���}#�v�S���A,���(�b��6y�T�[Pn.]�i��R˭���!$����^KJ�h��hv�|K�'A�Ep�'N�Z�A���Vuܘ·����v�\��b>�F���w��ߐP��<�b�}�F���O�+y��Đ;M~��M^k9%�̇�}c�������x_F�J3��Q�~��D�U��t�u�u�D�L�+�����A�[:@5��N�����I\g6���IⅭ�-A�ݽdU�K2�Bˣ}������L̴���N�\U��{�b�^�`��y��ů�Z[�$P�ⷾ������q��&�������9e;%R2#s_���(�3}�(�s��b�U���h�2�I>Ͷe�y�!�����>����9� ]�m<%�TD�5�� H.o����w�Ѿ`��KH�E&�VY��gI�1�=�]_ jGF��\S*����j&�m���ԇ:�݂m�/ �����Xw|�W&��}Ɛ^��c�ki�T:+��n����oj2΅�����D�GT�LF�d҂4�����[�����	�z�OQ�X*犪��|�'ҍ�V·��*|�}^2�A�6ǚ�tz2��L�6�J��p_�£�j�W�f!)�Y�a<������;3M@O^$��B��!�����5z��Tsr>Zu.D��d�Z�,�5Cz�I��
��Px�&�*���=�tϒw�3j(X�Bt��]^ 74��:>@�֙�{��|}�τgwX�����e�=vN�H�� S���0ٿ�)'�` ��2���S��7q1�x�ë��T�f��Hz)�ʠ�,��1�w��h	���B���J���e�>Gk�$+�����6�$�k�E�jbj����Λ����~J#���^G+4��JB(�K3�A�#<[��/������  �~)��f.��nm���$C���{�8�(��<Y:aIVo-1���۴�췩R֝~הd]��w�#oJ.�]x������r��m�t�_���&��#���-˷�t6ѭbPI�&c^�ш���ߍj8K�����r� I��DV[�oC�t����T%�vM\�
�{��a+iضa�Ѹ�b�O^��*�XeҵY(h��^{ދ�^���4f
n��6g�f^�
��6׿ꠡ���v�h�a�m�`�`�j'g��T�^kv�y<�j�Ӛ�����5B/��d�i�l���jO)��b�C<�VK����I��p �Vn^�}U
n�VNb1�+���<0l�l�w��bV����F�����9�&|�4E��9]�U��-���54wi���R�G�urQd��p��@�%�AI\"��4j�,\�w��-�l����K����B5�1C�B�.�^%�4��-��J��&_����=@C|�;�>��]GZ�5��L����b�OUݣ��}K��]���$#(/�������� ��؏���~s��\��p_�1'~�<Qb�Q��bv��K⪳�Ό��SD[#�Ժp�ž�i�"�9uO�0��Y�J������Iq�J��<��[�L@p����@����P�F	���ݰ���L���Z�w$�i�g ,?(���ڟ�{vCB����*jd)%�wN�G�X�3��u݅
����f{���'�1��D��E�|�c9>ɛ�r��m@5��Pz�%;D�,,�=F1�͔Cr�4��B��(.�j���x�_��F�5��{4#l��\�^�ۼ�P��XC��w�Tg?�&u���T�s��R(�A�P"O���Z�O�{vC�B}���Q.�I���цm7����2�
>�S�Z?�5on�D�b�Q�(F=�;X�f8�
��T��s=��u�;�Yx�:`�a��v�xk�&q�,��&X������u���I�������uG�6�	Î�04-�s*�-�p��@mJA�:F�����.#��Q.C"A-��X:�(z'V-~X@í6����z�#���n�to7^��~VG՚�K���)�`��˺����n�Kt�H��5w�L��թ���5^]{\F��ѻ�FG�W�P7_}�5&H"�gW�^�H"�_� ����Mu!����}�c�.NY��[ u�㪨˝���9)8M��)�h���!�B�,g��TQ�eB}JRk��4�Q�6�8�<oﱝ���l�f�'C�L�˴c��X�W �i������h�rX���à�\���T_��z���Na�O;�LP��h�{�����y��ҍ��y*9R��k���N��X�A�pj҅Z��s����b���umh��"̖j9�.���０���n�V�Z�5 GÕf�� �˅L���������H&]y!T=�w��%��fV�-�u:�@@Xu�\�(�w�>6M,D��I̓��Iv�M�*�K����Gum��UH>��/�S=�.c*~6/�k�~�>6�����[X*��s��T�ӎ�Dx�Uܧ4�v'Z��k��F��	FK����z4�Y�y��}[�����>#�ӆ�!}�&4��s���chH�\�W���0���[�Mq6��ɠ�+�uY)�P׭�8/��o��'��?�!����լ��i�\����:$.*[lg.,��kEY,��6��Z�ï��St�#�~�DF\��x�;�,��A�y�	�k�6��������@Zp4y�ݿͷr����K��������w/�<wu=-��jyKxԚ�%�gb��`��"L;A
�����4�Io���5��T.�49��~.Mƽ�C�d}SI�O i�ByL�y�4uy4cl��cH��^�D�r���h:{[��I�>����{��BH'�C����<�x�,9�r�
�;M�����0u��<��uu��4�¨�v�:+�M\��(.a�%;�C@̭&������$v�d�@�����XR�u�d����i:D����6.9���j{
�;���-hF�����3�!�n�	E�v���
�����*� ~�z��R����N�\Z>	!7wrl�E�?��%=�J��L��`ޜ��;�U;�x2�9&���~s�@�*�����D����Ɲ_�8XjfZחZ�W�I�lyo8`<��@&)��U�k8����R�>O,ų�Ib!O�_�<��BEȀ��}�p
AN����i�����d�g�ŧr�,�zLeÅ�H�%�u
�]�-�hmB��^#{Ĩ��A=��H����_�j3Β�9��dX��h����,!�7��Wzt��#�%����U�;�فM�*8�֚��������<�o?����s���N�#�v�<H�()�k�)��2�┼U{g���M<��0�xBWe["��=�w�%�jI�����^a��j9�G��(�-�y��6����Mћ�y���Qڀ�:�dǇ�w��X]��F։2��$� i�`��v�r�C��K4I���]=Ю��4I��&����#c7��������N΍�ۍ ��i�&A�/�3�	�F�Y�0.��./52	�������E
�}ű���V�]�)UuT�n��dIGŪ�F��S`����h�u���|B�ܕ,%L/�c���s�V���
n��Q<� �fJ�����
Q�em?в���W�&&4��o��B�d{���=e�'w�F4ޮ�����c�$>����i�/
"b,�z��0���s�o��-�ֱ������[�A��R�Ώ��qʊ��Y岄��T����R^$>�DH.`!�8�2bv��èn�`����P�H��S.nb�C��.v6%��O/(Y����q�i`n��u�l}��j��\�my-��l׵ ��į���F|k���_!�W��S525/��ҋ��rZ��i�� V׺d�YE���kҖ��5��3�SV��gu���Ub��_;$0��9$~O���E$��J����IVVz�׫呢c�	���� D��6B��{~�9.Q��|AqT��/"F��b��I\�����/�č&�XCR���/�\d��WH����R�=^-����QR U��ﾒ�On4�4����:����UA7[Ј��g�et�g�Ԙ��ks�A�-aB3�>�1y�uHMh��82�OĀc�Ur�{H�ql����Xh�Me_t���c���x����x-���s9ž�e�dE{�W{���L�������I
�%ۉ���]��1�%.6u����5�mBkA�J*yA'y�OZ�����ot�Z�U�C*�� ��:�f׊շ|�0���2ϳ|cF1�/ ���U����;[�����>ϛ�T�p�(����c�/��ցdm16�щ7"�����aރQ������#�ƄW��n!K�)BAYp\$���������9�Z�'�Zu���#��HS�Yi���~�Z�rN�^�SG�Rnj���$�e�ڝ���<��Rd��r.@~�4��V�	���LP!LX���6wkji�[���*!2Qaf�}��V�F�ٴ ���ʂ�'hJ���g]�\�C*�׷!�y���k-_y�`)xy0�p���(\�ʞ��7]/.��ڍE+N�iB�zbJ�e���r��^� .�׺5q���-J��]X΢��u|��{�6��q��]�׊G.?	�׈�=-�Dӎ�+�(%M��=�:?��~�h�XP����]�n)��`�eO�I�ĔbN}�* я�w���f��h���ZqA���"2.�=?}�\�N�����xe%{��?��/�����~n��D��F�f�>�a��l2����iC=޴�r*�䏶����В��J��R�ƚΒ�"�Z�{Z�a�Ä�#+�� Pv0��W �LWMx���dd,��?~Hr�*��DyZ]��	"�4p�}��yk��&�b��Lzߣ� �د��v���cE\}��^��u���3�e��̹��\�)n���2��Ws�5T��#�
��w�nF	g���5�_�z��ά����g
|w�go��f?���of%U-�%<�u8r��!D��=KM_��J�&���ܞ�=*P�Ykq�x���5r-=���1R�:�Y��Q�|�N<B����2�B3#��@�W8�p֛����7C�P#[M���Y���z}䚭{!�O���7D�.�����奺�|d:�Ɏp�հ�t��;��Q_y���sA�6�0�ip���NO�J��w0{������kV�ѾP����gLSn�}��$���%^����B|xN�����`�t�y�@5�	�k���(�xu_IΓ��Z1�"��vʫ�lؙr�j_P��v��l�z{:aݝ����S�qQ���@������ծr努=f��ȫ���Q;���(a#ys���7cPG>P1-=�l�š�A��ˡ����QǱߧ���'F�Ŀ�Z�X��a�@��u��HPT*ϊt�EkJb�zوt�E)���EW�Y���7�Sy��d�Xy� ���zH];�]�JC�{�zy$����y�9ah��Ћ�)x�<SpƎV!j��s��{�a��'���{�њ Q�X��ꁤQago��Al��\ ��$5%���ºw�/W�Q*��"�v9mtx�p� O�&��T+"�x"~�TnǼ.Umv�"D�O53�;Jmڐa�qT�X_q���=hJ��:r=�@������,�5z-�,ŎQB�3=�ؾ������bn��0DZ枂y�V���a'�62����c<��>�%*d�8�R~��^?n.�Q�F�?�5�|���V�f��	~r�`�W}�ٸ��u�����P��q�ފ����!d��&����Oyd
���	m��1�~��;��uX-�ɏB�[[���sn��\*���^A���\���;]���)�5Vd3��Tf�
�23���>�T9�8-o��-�(��w^�B��迲4���ۑ��'yi���GAC���&��0fG�}sJ�-v��r���:N�N�����{ca��i����׎ׄo�8=���B��'�.��5��6q��R��"�QP	�+�2˭���A�*_X�Jջ4�d���"YUƨ��0Ev�v�B�V�!~)H�I��s�N����df\x��B�]�A0>#�X�[�L9[<y�5	k,��l�SJm��1E�����#	�R8��K����&.�}-OҶq�;�DF���nS�dh�.+��U|U��p)C����n�tN��_�Ӷ�v�n����u`��#D8)u��7qރ���r�v}�v�s!��v'xJ���Ww��${��$n������s���a6�	��Է�s�*b��|O܏���;�}N��!/���>n(�im�ds�m�f�*�V�Њ-�E*j�53���n�◆gU�$,��*�� ������6�Z�A��������Fi�>�����1.3��J���*��I� !���|�]�,�l
�ݸo��u~��7��^�]|��r����x��Z�g�I'�11$��c���E �B݌�k%�d,��f2���g�}{�ΌJ)?��?�X>�=��.�D�"J<�L_����uI�m�/8�F��f4_0C�ޑ�_�c~���+���e\�ѵ�>j�aN�ڂ����u�����b
�Bru��.�`;�e��YIB� 6TEfH��+��/T��󙻨�p��C_�X����M��$����w@0�O'Ҕ<%�-A1�����[ AQ֘:}�贱�mX��}�-+k
?�:v#W�U�E5�@0��F�Y}/	9�3�RbA�h��1���"����(���<�e�,��$�g�I�1g�����]�´�*Dh�
=�wy	9k�o#��8����m�4a�H�������5'��
-T��5��Nqy��~x�I/��#:M�4��H����P��ka`�x�b�7�� w�>���r��J��>ە�<���N���)V�a��l����@� �4�nr��/��@45pV*t�S��OR}�=
��u�L�H�����y\�2����S��aH"� _K9��գ�+�B����V���S��`@�y�������9�#���[���w��<�?D-���%�^+w(D�.���@�R�������B�g �u�4�ʀ���b�G�z���&g��%��5�Ì�ׁ��[�8�7/l��iŋ['-����yR��.T=eH�H��	J h6F����	l�6�f�r8���YdʐL4W�|�[9��R	u��J����ζ�g9j����~����	u�(>�g�RP�k2B���WY���MX�~a����^o�[�~þ��_6n�D�,�jp�}���@A�HV*6���|���#�������Z�k]1Xb46N�z�U���d�/�\�3�.Y�p�P��O��ו\�$&Z'�!$�؏�,�1\���19�����}���WM*�	V�p[���=4y͛��c�Q�щϻi�@����a����MD���c�]�P�S�?8���+u��h88ޖ,��TI��]ĨGU{�H\JKܩYNi[��SBd�6ɒw���`:2��p�)G��6�{0l�� ������8
*�3\)]���)����ƃ�	-"�
�8W��}_�<z�<‱�ݺ�-�S�� '�=j�g�UPڸ�f��\�"y��s���Ev�����"���IaB��6���&��靫�AZ��V�r���"v�&1��d�RGb�E;� a�-��=����� ��W��������f��;�b��t�.��n���Ci$Ѹ�{�P�PL��r�3szd��֕�d=�#�*D���VU��@�n����̰���yR�=�[>M�ɫ~3�y�`TA�E~)Y��#��?�.BTvml�=ǡ.5��<��p���n7,eEMh��o�gZ�5�jR�%i���Y/�\��.9y1ۭ҂���2Ӷ(^%�T��R!��G���d=hS��\-�澿�v�Q�f��%&Ғ���Y#�/���+�U_�R�0;��V�>\j}�h�e��O.������ι|ǝ"�	��ґ��4���gF1�a��W���I�T���AO�٬5��dP�}�^�E����~:�,�1��e�2]a&(^��`a�ٻ�ۆh󑵚,�g�}��U�TDԤ���fW� \t(�PcUN��Q^]i����P�H�H_�}��U��|�M���r�J�j�8(�C)q
����Ag��{x8`|!w�!�-
���>���oD0W�'8�1�"�W�J��{�_;)r"G�[�X儸�z8�T���Ϯ
}3��n����*���o�3~����0�lUJ>e��|���ﭠ)_�H��4�νd<u^�����Fm���M���~�Xu!�m2��q攲}C���}A�����O������O����5>01�,���w�S�i{MmF\�Z�_3ȣ����w
��K)$BmO�eiĽ�׫�[�vZY�#Tv����R�Wi���򔟅������]��;�4y�����lQ�x��X�=��v^�=�is�q��9��^\(���d^�
/�V��F4BXtb
]A�=I�ΘN+h��z{%<�1**��I���<�XI��ou�\�R�|.�N�0L��=��q���:y�B#�!_��0��+ �-�ߘ�,�l�B��r�dIݟ���{U���n*K�g�|`�Ǔ�4��)�+���ĦC�rq�����
��n�i�'6�=U�<R�Z���4	:�2>���;������t���{�@��Qa��W⟸Xq�p�0|���5Q����CbE���`�� �����%3��X:�����},�*��|#h�CHi�2T�l�s?p�w��Lz�N��S�=y��q	p�3��B۩�]�1Q�d;J�Y'����O�|�>S�@}qm�mА�����J�g���7�ja�u�<�6)>�s\��XڞH�<�
�=����AJ��.�WHb���P|~�-�?���A�^�dz��#E3�ӊ��w��v7�Cf���6�1�����*��Y}�'\DIz�g	sj��;��8�c�|����X�Y��ٙ�F)d(�O��s=�ο;�٘Lժj0��'�Ɍ�@=|�g2'�M�4�jG�9
t���Y�C������_��8.聿~yR���_t�7eB3xί�$.{�Z�FѢ�˙V�[h+��$�deiB0�p�KƬ���Z��nv�V�/���쌳�z�%����>�y�g��Y|k�MqACf%H
=��C��ش�MN�m�O�%��wٞc"�٘���K��}R�Ob��	�R���R����K�\��# }���tժ���2��>���g��D=jlÅ�̇\��jqG��&�U�"��bS�����~;�V"��>u]�.F{�J��T����k1���@C����AN�xΨ�B�d7q����N�)茂V�?�م@#�梓Z�ZG�A�(�i�P�qh��9/(�Ŕ1��A���\��\f�fK3T.��<�x�i:}}��%l�R��J��OZ�p�~}�(h%�Z$Y�:p�RO�Ｋd��^^�rb��j.r�<����4��#Қ�/N~m0�_F��S���c�VJ͆"������������c�����m�@4;�5��C&Ӈs����f�T�4��O2دA�w0�Lo���2�ݔ �A��:�>��*�z6���˛%���4ĉ��ϟ�th2yR�m��B�߯��L��S�F�@L�w&ww<�B�2=����+p�lO}ʰ�I=���r�)�3/[���%�;zX��;�Q��]������?B��.��0 �]�'�ZS[g�4{e��x��i�[1��Btp����nu�err��|�sܢ��Јp�Il�������KM�L
�k�)���!��e&�eŴY\�' }O�ש+���,HM��`>E��ˀ 3۔>������V��E.�����h���=����~��Vx���{'�4�9�tU� �ܨ�D`H�7���pG6��<U��u�~�S䍭]*y��jA{~�v�R�����2���g-a�Z��%�K�^�,�	r0&��<[���[�H�J��~T�/E>���>�'G�&�_�.E�)˾'W����(���x���.b�s���Ԩ�9svXD�lu����!���oz������-�@\^��]�����́{C}^l ,�m�$f\^Z���n@]?�ǥ�i��=.���3���,a��R{s�w�&��ڞs<nV�R(!�B�U���;J��7�?�8�������i1/x�
%9`����u�~��).[W����x!��?��f�?w^N��<mc�zc�����Z���ҏ%D����'dA�G�:x��n�G/�����޲��wHZ��h�m�.!.����[#ƣB�:��JU�a!#��*�l[1_&��<�)�fwX�����ô`J��?���o4{�}  �o�_-�b+�������X��N�w�?�5(�b��+<�G����9.�C.��IQdz�^w��7V'e;%�*5|®ѷL�M��	�7����+-�n�U����4��+�T�� �d���#�^�咶}��b�O��˃����Z��,/�)�\Mv�b��AY'Ł��n��E�1��^yF��(pA��hq���m�㵺wJ �����!�!̑]Myg(ZK��U�G��H�=�W1D�ѝ�lQJO��jϳC6��Pi��b�K�VtVu�|<u`[�L�͈��ئL���κZrD���?k���Q.}�h��;����0t���Y�~jOW��dr��4��Ԏ{7����%i��&nO����p}�;X	W��Tg��t�x�4;!�����&甾DwW��OK�Ӝ�n��y����K�W7>�����
��"_���HPd�8Mm�5��G%��2ڝ�ċ���E��N��1J�07T(�l1��gwK���ĝ3��ϖd�+�0}Q�o��೮�߃L�ጯ�0�6�D�[s��~E �j������`�Z�F�z	Õ�e��_�hT��R]���jU�^#:d��΋�Z��9����P����q}������_�cN��D�Z�j���9woO�xz.�c,�QL�qd�-�v�X��D�N�f/@)9�E����S�`D;�`��uwx����������K�P�"x��NPY���]HA �,�M|z���H8�*w��ɶ|ݫE�9,LYAۿ�x@9}�sǾ,r^��w����]���G��X>b�$���P�8���{AkҰ�~� m~�`��Iԓ�5`�Itp�<�L� ``?����l!	*��e�-�O�����x)'y�Ԑ�9��@:�cpE�'�RY ��ܙ��¿��0 &�.�&����w�m�qAď�,���ם��̞��݀�R ��m�����ꤰ1�vy���C��>�G�K+�X�,�Ր��$�/���9���)������m��N��P�x%����U��jӤM+����˔|_����K�n,m�
D�,�x�˴�&{�|jͿm��2��h�2���D�"�+��ߡǔV,���kc�ܓ�l��?C.#R0�:,R���� J�o�J��Q*�r'C�p��GYyA����X~�FT������'U(���;���>���Pc���G�/'�Sb̼Ӱ�@ y�8�����1�}kz����wo	�g7��^�L���pt0ݍ��9%<M�o�%$�	?�v���u>}Z`�ov1��enʑW/����JC ґ�Z�c <�ج-\Ok���h2ӋFz���ij?��c����;��h�V��7�7��e�˫�f�!�\h�mY�Es~���3��y��YW�EBPމ��*
p����Y������들ڠ��M`K�7�=*��8������Q�L�͈f�����=����q�]���w� (Jw���x�1�9�` �4u��+�����#9��������]�c�>ebU��ڌ�y�����`��yB�y�T�oU�!j$���_�&���DB����_��C�=������Q1Ô$1g��9f!0N�Q��G0T�Tl49����[��D^w��{�)��v}d�;�ZFSO��$&��/8z�#�zÂ��TK_c��E��э�pɍT����y��B+b��Ъ�?e���>|L�z�^�?�o�Dv�3��[���}���$��0���W\�S��?�������;�Q�V<���l�F���B�g�{ �ȿahw�l렯G�y=v"��8	�>k|����S!�N�����;����쌫��9A&�oL��23��yz������N@�?5���:"*��`I�� S�T_e�,�ܧ��*��k�S�X��\&+��R��e��+<�MÛ����q� s%t�J�vU����~�.D?�aj�t~3�xأ�l�X����i��N<-�Ԩ������69W��!I�j'++���"�q|��TB5r�6B�A���"��R4�<���%_r��#����Sع&K>ߞ&a~�V��Ȓm�������"p�q�uNٛ:�����mÕB�Ú'�m"^n�?�b�TQ�R�k~茻��!����Z�ޠu��n�
�r�B�&K٪{��@�~�7��*^�N�LjN͝�Xm;�|�����*S��Bנ�7&EltE�4���33F�����6M��`��\�W�K^�Ļ7q�:{q�~��ˣ�j'O�G�63���$��F��5^�������r}�I�?.�R��%�X�k�}��b)s���hIm��C��tu	A�: \�q��Y��9�>��3�2�O9E��I�-�CN�t���8����v�0�ڴ>�����{��z�B�h�x���2�����w;𼋊+���2���m���hb����E���r�����[0u�J����v�GwrD:ZT2���J�=����<��+>�#���i�״إ��71`&�m�MP/�V�H�`$"^D.����;�"Jߘ�UC�:�X7�|��-���zm_:��Fb��!)���)����v�#e�k�����EfYhu��`m�[�������8	;����-g�SBHen���>�|���R|-:?,yc�[
!Uæ������9�,c9S���
����!����ttmN?q��c�Rr���e�����D���?��x��~��}������)�\��H�����\�F�J6� �E���E!�f�gp�h�ԷL��f���ZG���G��'�0�	NZ��bOE,��(G�P�,�L!�裱��o�
a<�!��=\fҧ,%>ӻf��j��������6S�a�e��/ׯ����������.̯v�3O��nl5|,%Y�����;�o��ᄼt�U�R���r(ו�}��C�ڢ\�j��$E껸⫉��8"@*���=�Y���S�#��Q��kfo_�i��)�9J��A��Ԛ�m/)w�>�p���h��@,�~)�3���u~�'�1�����lX&]w�22�n�|�^�k���4�����ۥ-�N�H�m��\Q�P��-�k�J��'u���א?+G:p<)I�t�w
sl��
�[��(��u�����	f�>�%�E,���!9��F=r%K�M x�N�6�̆6ǝ�θ���4ކRsüm�����`y��k�|�beP�h�<$����YM>��$��!47cd�=�R��������6�]�����z�z��*|�=Je��m��B�C��8Agt�kS�x��){�R_],���BD�_�b�r�Y~S���YlI��n:�?2��H$*�����	�A	Q�a��A�'�4�U(��F;�?ݣf;�
�K�I|�'�N���Z<�V�j�2��~��^~5޵L�6c5�Sj!�ېxT�_���z��S:�7�*��x��ʚ���[u��Q��va���͔����l�T��!��|�eE��F\�gX����T�&f�D��ɞn��E��g�ԙ��&�J������}�B�!Tuc�flK�@�v)��`���CL@��b�Y�y����/���<Y{|n���m�kȄ�(�w¼*x>�,�"��po5�Ga}��΢V
�آ�h��:DK���wb����lK������pJ�j��-�F;��iF����[���K�Y�6ӵ�p����� e�+��A@����ۀ��>W��X�m|kBݓ&��#��W�X�Y���������	�,��o'mni�Fq� ��lOԔ7�]!�Opy��J$����]���RDzʇLq�8 �E��:�~=B%����V�oۆ7(���WAC� ٘ڐ�L��0�m6����������'K<��eͷ��0p�'�^�{�{�6�8F��8��3Ȉ�N 4]9��!�.�Zcƫ�<�s�d"��Z�?2�4��D�QHt�hU�K���[�ȓ����g�ō�[���\|��5��� E[�MN��:�I\������Q`�-��mHY3��\�<�����'��Jv�%^PZ�j�j �=��vD��S"
M��%��p�~Uv���!�)j���z�mV�1=	�w��X��i�asLY�2֐�F�W����N�J/��2�x�1�>nʴ�:P����fir/�?lf ��J#N7��@��ރ�$މ�dS:�y��"aް�߰�<6�vĝ��D/lv�^}7�N�R\��4�-Z=�T�>;p_��/L��/@���z6�X`i�`i�.L�P)P�iW3�j� ��-�3���W��[��F 8EC���z�,���Tޅ`r[Y[�ө�[bz*�d↿�%L�zlb�`5����k�I*�j��@6K�&둗n�d3X��}����^�0%���x�q���k�"�䟤ܥ��S���0(K���	��lk�C��}'��e�ׂ�"������y���L��NbX�ie�8��`%��]�]�|@��,�%�֟
����,*��5���B�6_)92&F͘��X��n���m��N��,BU0�¿͑�7�{05p�������,�8Ṡ'xB[�F�����Pt[�993�F�X�����	�Z���s�3�L����f���Z2>&��sqs����6��<W�B>ǩjƶ�~e��l8�Qt7�/��t5 �ܱM����4/%u�X�y��z�ݫ��jZ�l���W/��/$�`2�|�b�o;~�v��Rݹs��2�Q��K�)�֖��d\H�xP�5$ᱼK�_ޛH����2��mhܿ=�c�P=�+}S��I�5�lE����'���{$�b2xej�ۺ���������,���}�-Y)�K�������s��8�܊��q�ox�xrjmb�W�0�(�q�.��h/h�"��떍�8�<�X|�7���ºK�1'a���Ǝ�o*�VE,uAOco�q�>�4��>¯S��o��C�m�0ct��q	Ѫ����}&-I�WQL>�pD�T�PU(2r�꾬PJFU��/��O�Z{hvC�W�P,l�6s�
Ww��4�n�̴�8͠��=,'����x�8��؟D=L��y{���I�P��b�Uwu��	���^Xp$��Is�B�f���)�Rjs��Ul ��
�3�u�nR��� �"�֥�ìM_�Y�[W��(�*
�{{AyP��������������.��؝���
s�gD�Z����~���hٕr�9����ќ~M+p>�IѨrZz�;��>��!���゘� ��IUKs��Ta�26=W�
�ﻣ�DZ�&ƹ���K��8�"s��E�S����QTN��:7u�J`/�d�p�8��f��O�	���;�q�&�ɻj2���(��%N]R[d/,0��(#.�^���{�΍;P���/U�����:��Q"��� ��PGߠ��j�x�S�ـ����������|�����UE��Eㆧm�Q�(�޻�a�$�6��/�*�.���u��j���IɂO���f�\��V�3����>�'oU~j����_t��.�:��v�A��������@�L_b��[�m�\�^q&��ͧPC�P	ng!��A5�@��ӫ��6�SpiU��
j����\�Rַ����>�fe%2�|ٜ	�e[�i]��H2E����<�P�|z~fQ�AQ4=�2xťFK����d�"�bo&��k�:@�P_��|�G�1\�h+���V����9+�#����i����%r�X!7� _4fBȉ���~MS�����gP��}�6����IAf�p��h+b��q(�a4��JĮ����6� J��q��A���6W��\���:�3 ��(n+F���|4Q�/k3x�d���Ğ������?�L-K�_L��qm��_�x̸} ��듰��Vg�
�%3�r��z}X�*��y��G���V�e9Z�n_v�eW�7��nϩ?"��N�CRl�L�LúK_�U�K��@�zL����c ]p[L�EubF�m���&q�.p�-B��@�%X���bRF�F��>� �Or��0�S.�%<[BO"�YE���lUp�P�v0D�J�hs!��w,[��1����,OعmM�&ㆵ����ހ+&�A�s�Ks��Aa���$����3������m��'�Y���+�)5�-]�ͪ�:��^���ѥ�x��F��ܞ�J�Q�D/��jt,ֻ'�x�0��b���R�Ƒ�����]j���|� \���HbO����&��ۃ����H;y�~	q��eO���c-0A{
5�۸?}D)�=�(%h�P���k!��J_���{�/�^�n�$W�D�����1|�_P[�f�͐��*@����s �
��h����!͵�m]��c��9'73g���dSG5y2�]���d.b�I?y%#�VV+���UB:�+>��� ȃa�@qz8֙y%��<����޳� _���;�FT�s]���W{/CZ*4����Xs\��U�"�B���
䶜��`u�X3��$f������"�<qv��3,���K�B<�å�ǹ����OՃ�H���q��#�C�u�E2�X2�@�D��c	� �DD����?/!�5rA������-nK�
������g{"d�!x~�X<��5+6zh����j��]��W�������A�zjZ�ge���#��|���+���� �_Z *�L�����5��=�dN�6��m��=��v"k��r�P'a*q����8"�kͲ]�#�3��,�72�%�(X���m�k��R*fV%�w�����wg���4M�;[C�g��-�o�9Z�I+i����	qo�
0|����/6��$f����CE��'l���h*a	*9��[�W�LS�74իL�*���O���2!WZ2���D� G%X�Q��c�71m%��[#}T0��_��A�Y][��l���.��\���M��=��O	x�%XK��w��Y��Cȣ5u_��bU������)��*���z���h与��Zѧ��]���`�[�cȅHck���l�����x�疐S#�cƼ$o�z8��@Z��ԉX�U��<ƶS�}��L�oOHq>(yrR�d���&P^[(o^(l!rV1��|}c$�p�J��}dK�����y!���m˺��bS��:�Xi��%W|�1�Q�����	���o!qRq�Z� ^/��`��=~�{HN7��֫m��X��kM����Zb!��#�_"�����PIc�N�vF���Y�m��qZ�@Hmϥ�%��O�<,�0b/��n�w7i��f�	k+W(��F\[�tq�3:�e��ޯ[ܣ�V�إ�(n@M2���ʂ??�}Ph�S�p�f��r��,��Huݠc=J6&�ÕO��Blx(�r�ɕ���̩�wʌM����î���k�n�pA% �.*���iTïu2M���<+�+WO⻫����߹���1V֒��#�Lʠ>�pa���7�2����T�y��5��S�,�Nm�]�ħ�����F�55���NF��/~��s�������������,��U�%�uղ�~�S6|�ꐥ�`-�<y
x��
t�>g�:}��jU��(�.�aQɤDUѹ��f�+4��l2����ׂ��*&K�����i���YK�p����7vF65zY�k�� ԙ��d�5 K��kM����D��T�n�'��|���A��Y�A��!�f�X&ع�=�`�OD��V�@3�SW�{fJ�&�nҹI� ��kj׊�y�ç�KwY�ZA���pPw9�U�S�
�a�K �S�++etnXzG}SN47��(�$��7���J���E"��W>ȁ�@���_�RQ�ad�8�X���������<c���"x��QO�z�A�yv��������Q
nrG��O�����o������[����, �^�X�|l���E'�4F��B_�t_>�����^�_q�G���q7 ����2�����rI�!���4k��D'�c��?�����x�H�$7�Ҙ��������*����"�p�y�oߎ��?�9��{�P|�$)�K����F9��9~1��w1�+�P��m�F���U�#����z�=�r���];���m:���@q��	�$��E��x�Y,>{��Y�g���5GB���	��娧7 �����,��\"~���z{O������c����t�/4_�z��S�4&��m_ф
�1�u���񄢨H�딳a���o?&%'�,���S�;�����6]� ���$On�dѸ�Ȕ����٩�ܘ������Gy��_�e�[&<JКB��%G;��}p��^2������@�"�˕��^>��=�AN�ǳFI��g�/�H������l#=?&T%d'>Y,���T�圢��GqK���D�vջ�u,UamRF�Z�m��nE�_z�+���:��˯C�MY����]md���8�����9��f�����'��/e�H�'�Q,�tv�Qg����8���>�0:�i�נ��)l'6�d�3�Y�˭n��"?~�Ⱥ�H�P������x�ٖ嬖��-Տ��9h�v;�	�5a��ظ�ssS�i��Q�?�J}ni@M4??n�ћ����381-H8�'\�P��#`�]�8�[W���F� i��Ј0w
�����~�e=�r��Bɳ���T�Wb�K���
�yx�>�[rd�p�o�O-3|���4����rW�v,SS�X����@S��M��:�V�# �,��׶3L��8���%i�ƞ�u6kX �����^��[�(�y~�0S�_��Jr�~1�P/_�I/�Xo��)S�����B=$��^BH/!��bD�3hb�[^S?��ashN�O����Ⱥ@,bV���=�1�崤yn=���E���%;F��p_Xl ����r�����٥d+�/���V��k�;E��e;M&�	D����C��Ti�nx@�n�;t�14���5�}ަ�֗�n�J�'�kT�˟Ϋ>횋&�;�}�lS���{���z)lEX�w�d�*����y����-��N=$����4���P�]ʗy6���۲�|�[���\O�t�[��J�igr��o����zk���&�ɸ������M�Zڄ���XFr����4�8}�}5�֜d��㝚����N�ןq�{�� 65+��;ABH��1�WS*����Pky��Y�xĨ$r�P�_�7���l������U&f��z]���P�c��}��h����;Uw!��@Y	6��&���˶�4,�oVE;\҇��%t�`T��41�W�*��4'�c��-Ԯ=�4Oڎ�f�����!��������+�� J�i����p�-ؒ������:7e$w�*�7y��$�5��T߸���ء�-ߏf��mz���j[q�Tsy���&�9�F�	�J|��SZ��D�ZV�Vn��
a���BI�Ϡ$�}t��k�5j�$-�5<]�x�Hp���]���1�i��#UsB��D*g`gaR��X!H��[������Уfj�P֡��n��<��Ʊ��^]i���"�O_Z����U��!>xx�*�,����*&�=MԀ�8��EH�]a�6�hp��e
��I�TG)t��Ĝ:���%��7$�=��Iv�n�����){���˸�`5:�?M����L1V���3w#\����0у웸3FgU�	��d��FC����8o���.�	]=��G�?Ț�Ͼ5n�!��,E|j8�ŧm��Q��Q�B{���-��`��^�ΐ$�=> V�����>�	��n~e�4��܌(5ׁ��=p�� ��љ�ч���7
�$F�[��p�BwC�=gF�{�.���q��|Ο@ȸoT�"�@$:�ߏ��/�����e�����N1{��WП��Q� l�v��wyZ55����3��}��#t�_�?��r\�+q�{c��y�ӳ��E���h#`��í2)$	z�,u���y$�r�XzT��t�3�~�ȅiy��C���4�w^�EEf6��i%iG����OY���.�������#����?����l���pk^[�.��_Wǈ�� 5�2�?^`{h�Xzq0��GؐKV���]x�3��~K����֨ɕGA6q����Lkdt)3!^~dן��T��X�f����2�)ZQ��胠�?�WC-'��8�I�|(� �`c#�m�2e���Vf7̦��bwc,7"���%�*����5G>���)�Z�J�+,u���Q�'<�����W�ĴQl��	&b��Pfp�}l����>ʧskX���#K`.f�r�o�O�����N$�.v@<�3��Uy���(��ܕ��D�3��g��pt����B��{u&ˉֽ����ϱS;�����LL;�V$�[��ߊ�{}�Џ|8ǩP}�L�Y)>�[�6�x`�~Y��"?��s�AѼ7�tS6�b�� "��/�>�ě"?,:��23�˿���}�|-��\��f4�3R�:�<b��ON������Yب���M��7��3lL �CN�G�X�Qi�#�ҫ*�"-�_S0ÇU��آ?�s����NQ.wF�+��f���w�K\��_J^�3�x�2�������:�̩��[ҿoI�����Oq�~͒��0_���xW~ K��j� 2ˁ���|/���Z�sw@��E�VΨ�`��t|�)K&�0��`��Rq��n	��f��K� �(��c�.2�(�@�j(�� s o��b,g������bp� �����)}t�p��8ej�jw{>�f�wu�#�*�VHΆ�;��Yا��9�W[�p8zf=*^���c�� �T�<oՖ��8��_ަ�<��!���K��_�kG��3N�8��*�Sc��.<���@�Pj�H(��(�AL�j��.I}7kd����HCp��ȸg�▆XW c�җ��H_�6�ޖ��|z$��K�FX������,P�0n5=;�j���T��
��uC��%�@�}������Ƕ<.����<5�D>�е���rt�v}l���R�?�p,��:�r��1�;�/j��כX���2�E�ћ�"*����
�K l����d����½�[t~�:�nQ2�Ờ�_3ao�e%�.��[�K��Ͻ�r�."��Tw��qj�c����Xu�n����fF��jį�y�n}Fc�z=�hF�T����pvZ��Ȭ��G�紮K8B�f�@�jaVIVA� �pk/,D��t��\�_��}L^?m��8c�P�N�����Q9Cm��Ű���R[��n��B�Ω[�����a��' E�`.�L$�Ֆ������:=�����Z��EY����ݜ\ޏ��QSLZ�'�Z��Q%�ܞ!����g�z!b�D��"���$�*��|�0��Ǥ�ſ�׮>��x�,���cb��g2lz#�������t�)�����I8��mi�����������gNx��j��&�od��U�S��έ:Ҹ��u���>d��yߠsq�Ah6q?N�K�j�����f�`v�ָZl�~#�?�s�)��4��wT�O��ͷ�M����ŧ����sC3�"lԝ���ݙ��{��>o��0��)�������2d'��^�k\�����j�ݤ�kU����Xq,wg��B6B��������|��ECU����9ˎ�8�T��6�\�����4��Z}�9����3e���2�dm��f�I��r�/�C����X���:�YOcG�̳�l���du˓ �J���=�g2Ur5Z�)o0����dQ�u�k��S�!m7�m�3*���/�g\9svaZ��������]3m~2V�z�lV�tL0'�eֲ�å;V���.�W�㈟M#�9�ץH��#C"aG�u�R�Q{VL�
�!='��vrDbl�Nt�		�&v�X�`�s��9�7�u��wA�h����2��n�PT�_nEƼ7\dh���<��O����[q�3Oa]�{�Շea1Bb|��}���Z��i$�I�C�!�=��5��	!41�p��\��L&)n����tœ(ַ�K�P�1���yGP�e�x���p��5�ز�T�+}����q���H}����=��U�����x{�D,5A���0�Y%�1i�LI|U�K��tK��y+kq�\.��q���F�wL�8 c��ğ����}����t�jk,D��%�Bs�^�ơ5�����%��=��
�� Y�7�FN/'<F��]u���P���\���j�n'Nٽ��\P~@$��Y�wẗ́�eW(;�$��6���*]��H�6���P�n*��X��Y����3�-�Db�a�)���&�I�������x����l�s�����}9ϴ�,k�K�T��Ӂ�A:�Ǿ��ن���&+`c���q���Ee���5�7O#� �%�ƶ9D��^��?��(t�j��D�d�Pe���Oh�`lT��G�>2^�ԛ�^śK(�0����*X�pgVoC`jd6a�zS�X�^���8G������f���蝹��,�����K��b�{�z�D1B�o�0�.k鼹�e����&�~� Ӥpy\6�=�A[���<r��ˈ͔w!|�CC%����˹�e�Wc�J��5��	��X�[�H��vs���{=k�;�SgU7�hH}t��܈���@�{�pBX���f�������cB�Y�)�l�Q��4�ھr0xV�P�v���K�����h�{���]�������Z\�*�ߕ�c1�;�AY���3^�>̉]���ꈥ�L����}��H�>���kb2	�5����%`�SZZ'�V�0���﷡vJ��Ѕے I���Ɔq�$��вuXu��]�q;g�]��ɝ�Ԏ.7��ȳ\���r�U�r4y��T��o���"RNH�O�u�Y�]���Vl<��S��̀�)(-Kd���6%�W�VŴZ����VL0Z'6�w��B����p{�m�F�깈jY�$ܮ�nڹ�����@�$.Z�U8u���j�{�4��8e ���~B�o�}w��؝-���y5��}����[YzDs	3]ݬ)ƣ'��T$�f��O�Q<�w}V#�����\�{ NqQ<4�I�<��jP��G"� >��iY%�oE�5fV��Aox���M�\��5Kxee�OU���q�̠&�|2N��p�M�:U����Ԙ����R���z�1E�ѻ�;G w ɖzxS�kj#
�3�\��)x/LhC�F�YǸ�$�"��?�үO�rn �O��0�_�yk.�G!	_sF��8�Y^��<R��̂�I:L:���ԖP�ɰHJ����)l�c�}��N �������h �v�>�t�tTz��:��<��H�u��P���V��r%����=��?n���ǔ���u�0���V��K�Qxv|�'s����w�\lp�ZB,�i��e�N�����%ҹ0 ��[�e�ݡ?s��\x
��g��b���h��I�Ț����[XM��~�k�
$Y'���Sɍ�U�.���ս���]&n�h���}�6k�(6���<%N	�p��s�*
m�)qV��\a�i�����$�M5�X��]�/5���\��xg/@̂3�Jh�VZ�n�JH�u��şK����]�:�!?+j�+x(͓�mu��3��Ma~MG�
.�TP
�$�,4'�_�hi�륍�B(�k��n&��1�����d��%���>)'TBF��v�U�t�)�����s�W��s?�m�כ���4��N%lX�1�dO\����!��|jymz����T�,�]T�K��ƨ���*����}�h���&��J�s��-�W}g�j\݀�v�0g�]�mѡ�9Z'ԏP�ȮR/����X������m"�C}����9�B�lL������95Vvj�(]�j��,�H���d�+|4��+I�V���,�F�~��q��,���U'��^��[��t˔�+i(P���ɃA�W��X:Qm�E�e�&��;4��PhV���3KH[�r	�Oy����l�����y\3v�����<�����s?K��t�Ţ�Q�l��	¡�����"�0��vIaI��菨j^-p`*C�UM��e���6B%D�y�W��d���{E� `�"_וE�+�o���s�fE|Xf梻�Q�ߤ�ԹPb��U�e�SAU~�<ݴ�+Ih.|����w�6R.^)�G��.�AT�4�=�����WP�Yl@2��5�v
���g��'���%:(�=����s��j6	�����-�\~li�}���ՖaY�A_���m�y4˹v"8w�c������_���YD�I�0�mӲ�q*v������3�<<n�	���G������O�j.ɪ3�w���	�}�EyZD���Hfa1{ZG�㓸<r��.���*Q��\�yfyq,C��b�腙���h��d�A�E����@��b3��؂љ?	��	�!2y<bÓd��ҖSs)α^D����em^�4,q�)ȉD1���u5��trV,˲,mD���f�mW1:��P���ס���D��"�S�~} �Tx+�n�ɘu06�c�qm�_8ƣ���,,���G=()\"�����P�&���Ƭs�k�a&�$`�it��x%��� �9g 9�ñ�/2��\�B�����4�s1�Wv��^�{ښh�r)���\Ԡ�Æ�Ab��Wa�7�ȷ�X�>���!_v�Lq�+�Kx&��֎h�=�F�tX
�d� �,@����̼��Ņ�!�ҠZw��d��ِ�3梖�>�[<#��@�B�*����/��{��t�~�9���k`�f����&%us��6T�0}�!@�v`	}�/��-�G��
���7y����-T��,��6\yZ׷^�8;HH�/C�xjX�pj�+I1ĉ�8_rk��<�?�Ś}�4�aF\^��h�����@s���;}C�2���j��r+C?��u�q�ŪNG(^���Fi�|�黻��1@ZE�r	��eN�*K��R�N�%ֶ���q�j�"�t�����Ć`N%U�S���w�I}R�y�+�(S��c����0��e ?�֗���� ��;>��l��*�n��>M
�t"d�7��2pz�=�-��I��/Y���*����ە;XS�)�jh]��A++�����g�aS�9+����ŭO^������k��Ab�j폕�#��bE%�N�:E���2�,�7u!��=�\��"�c;D}C?3��j�소����3�S������e{�o �1���ɝ�8�)Uj��$�g���wI���Lu�q�����ÿC?VV�S��u 6CȂ���Rh��I4�, ���I�x0Q��˔�^�0�����4�1�$h��f��=g�"�U�O,8Y�����)������G�=���LF5_7*"/KB��=�Б%�����{�rq��k�ⶫp_�C�¬5��p,��_Y&�֙�m�DT�R+FA�gm�H�?�ŉz������6u��}ܑ�p�S��)��~ X����"�R"o�������!��ST�s��J�Vxl*|U�s��?�Dd�8H�G��/^��j���̸�^����>�Y��\fX������&7�S�=[��]n��Њ��@�����D���ҭ-O�v0DƵ���Ú���Tˏ@�2ݧ�Ѩ˺����OŔ�+���u�rq�,2��"�%Nm�o���O~oep0H�v�7k���ъ2�Ka��+�J�T~s6�a%�bTP�{�l�(�/�J�<�AR�e3%�� Lrν�ԁ�z~�ݒeY�j����*zR	\7%37d���t#�c�'}CϿ�)�ح2>�~:-k��v�?��Z�n��Y�$PZ�b���&��]Y�"��k:l��B�#\�g+��Ln"�B�]TsN�C�l1�S�n&�c��|vk����?�qm�߂Z͘w��`���.�4P�/�Cu~�o���yz�'�������N� F�y�;��Ӗy"�\d���9�5��U��C �icI\a˵�m"Eb����x�2d �[qx���\5n��GH��l���`Q�A�
}�X����X��[�Dȡ��t��E
��$�0"������=_OI�'$��K�0pT&��n��6'P^rM�˳@+Q1F�x$�c��Y����Z�nB&/�&}���N? �j<E}��[K�]8ܥ��$��Ψ\gFt2�^����1���ު��3�'�����5sj�÷d����r!4u�/��!��FT.?(��K�u.)�Q
_h(��$_#^X��B�1'���D'm.��nM����z�5�?;�K�?��;�<1�[-�m�]�a{��^-���q������UH��}$�FF�ſF�������ntHK�V�'�G�e�2B;���M�Dk��)�X��?�k����eu'S�} ������d�_!t���Mn�:��|Vw��4�eؠ.l-פ�$D�rUi	a� ��&[b;0�s��Էޏj
�E1�̋U�uy�\��+O �¬�A��A�9j,P�!#0��ƛ�7����p��M;������ �N������D���B5x�<Jjִv�p�O���?V�0�_;����)�~��n����J�5��52\�u��uo����*_b#V6z
�j�`f����ll�.�v����$�k�I>�j}�C=��r,c8' w�UR��s��K�	n���G�63e��t����v)�h&�G��=^I=�$e8b�wh�Q��$�#���rv����'i~�R�K�Y]���) �\��K�ٽ���Ow�o���)ʝ�Cr���
m�HTjy4�2�g:hU��ͅ�����W�h@����	5��( t
¼tN��3db_av}��&�9x����j�����10
��Wh�:��t��ѣƑ�#�P�_��gg1�ϝ�X���9q�;r�5P`wC}����L�J�1q�%��1wm��F��{����{���s?݈��,��}ٲ�$�bg���I���89�~70Z���Q�����(-g�*��^&�5Mk�˫�+�.Q+Q ���XS���c�v��Xh_�O�X����e�wΆbG�DS�犃��3��xӉ�����*�_5�z�w�p���uqLZ9�xZR�֕j���o)^>6��ǔ��Eb���P�:��+��[/h�C��n��1�ۄ� rY2Z�^y꧗�M�\>Xt�)�B��C49h���/�y��NwA�|���Q��v�WF�$��������[��`s��X:���B!DXW�o�RQd�6��l01�.ݟy|ļ�K7��
���N��zJ�Ç����E}��:�1�=��<33��6X���6A���՟�0�5�+
]�e�|���%B�.?�C.��G�5u�ʲ>�P�= d.��QVa�^�e��(M7�S# ��P۟
1��R&k��&���V� ���2�n6��1N9��Scзc��	{�1Rͧ(P�	R�)�+�����|�����w�ѵ�j|��"f.�[���	o�F�2��r�s-��9t�~���E���5���=�
Ƌ�����*x9A'6����p���5o�#�!����6�4��\��icb�!��q��n�GIu����e
T��=ց[�J��eͼ]����7e
�U
z���Pb�%Ũ�yI��+�ș�jȬ���@_rы�m���<�yxxu�w��p�Mv�s�w�����}]֛�N?�Ee�;2���XŬ9?����dT����n�����G|{+�@���B�mZ=:����D�U6��FQ���~�2�1��O T����K���a���5����9� �{�U�(��ؖ����6�Z垺���.nW���K��!��(ӏ����������V�1Ґh�5;�/ۇ��1�B�M��S��͖�#>P}�����9#FCeg�>W��Zf�s$B�`� �Ø�����W:�캐�e��:R�Z<��Ui��	B.+����:<�6�Ȍ3IR��7矵�x?�V���HQ=T�� ��ׄA:6���}��z��~p����>����m����@�f�>��Q���V�">��H''�:U2J�߆�5�`|��L"<��w���>��Q1���zòy�T��K����������B�Y��}B���ݍ	W�M�@|:J���_����9q������jg�/�^��|N���0L�W_$�~�V G�iy  �����O�mn��,������9���Ŝ2���^��d8�%��OX�v��2�큢p��$�����+k#OS��7��,�z��H#��3q��gsx��
F�	S��:�=�+H92�8Ը_�w�ʻ��dkS����?����GE�(�cF7�vh~��K�y���dG�K���c�%��VՎ�;�Ҟ�p�Q9#�ګ�[e�?}��`�N�E(���B^�JU+�"f�#]%�;��x��v2�B/y%�����D�sF���w��d�w$���b���2�=ʏVWi>����:W�i�^�߽���c�쐤�'�j�Pd7Ƌ���h��^�+�:&��tf���Oy��ZW�w����$8pp̀�d%����O�U�������oB����}����.t4;�h[��\�Q����ȭ�EXs)�ߘ'���Q$FE�M���hq�D�j�1��g��1�m	C�l�qi^��Ø��\� �??���+O�j��� �	�j����˰+4]4����z��)���^�a���­3q{�}[1`.�8Ձ	�����O@)m(f���-	^���s�0�'L)�� �wpBN�</]3i �r|&`3����-�Fh�^���6w�i�X�����N���}��6��O]��ފ���*��ܺB��&g�� �TOV����V�Fjd*mԁPe/?S�z����T`�&odl�ڴ*�}�*�:2��D!����z�9���/�����:Ϩ;+�(����-_�t�`�ydQ�d�����2��zD(NB��q�����>�u�H@�}lf	�a-����9�d)�,�
�ϑWBz�s�ܐ��Fp��K
!~A��/ ~�Q~ܳ��a	�2��v���{����ЂM���.�9-� ��R�P&���T�nN���y�eQ7�~(��K���x���'�\k	�(EV>i�� Ż���v���"���!Y��+<�u�H��z����xA �=��.|z�-a�P�옥x&!}�?�\>�L�V��'eK{����U7�#����И,e��a�M�FT(%3�aY���j�4M1����W��m[.���f�F7�Ov*Y�92kDo_�2;3��̠��"����PQ�U���_S���~/��,5@Vq�@&W����n�L>�����W{��N�\b�BN\��ީN�?M����k�|9A
�q]�n���9B��bw&��A����T-8��t�ғ�G��˺�Z�����Bd!K*.Q��r���W�m3�T'���6rHnW�u�n?;���Oe�䨷!�������]%�Iz�4G�l�;d���O�,����V�:�\�6�Iy�ߩ&�i�!�����dO��#�?�P�j�ў��jQ�)&�?�%q�࿥���7c�w�@!w�Z�e�}���I��\�kR���E�x?0������_zZcw枯KQ_�:�uH�Z���*aIc̈�p
��F�srS��?B�� ȏ~���~0IH���7H]����9����J)�:�"����G#��j�"���h!�!7�'��nlͲҶ$<�v!���@���i�aH ���dudl�t~�>��&36Vd�� {��X�lّ^)��a�ę���&���w�oo�@�������6��[sp
O�J��~yL�{��� �Є����f� �e�m?¤�|-���ƾ�$��J}.�����p0�3���H����ӣ55y�4D�6���GR��h���x�S�E!ƹ��~$!/�~Q7�]B{�����F���2������	��0��v�"'�+�m��%c$;���Yn����T������f���?�%ьX�K�8ϬH�-o�nr�]�Ny�r�oˎ�����f��6'�)����&a���T"z[���]�������j��S8��t����J��fuK�tev���e�C�MD9���:�RA5.� #n`R�%���'jx��4t�Q��N�[;!f�-��v$���#�J����J�բc����w��P���٘�a\��<?j��KpO��D��6G�����G־;�Ϝ�7�m���C�m$@����� Ó+��{�����Ӝ�#��:�)VR=�x�ݞp({Y��{�r��8Mvv����������伳(�]���3go�����c#%���S/��mI�~�j	�@�	���=�'Z�!Ђ������,�0U�09�[��g�%�8�<��$���Oƞ��dD��+o����H����G�I����aZ���RKxx���m���Re6��3?�_hm����L��ۃcu�E�E8�����X����0sR���K��J����k~�[A4H%�lA��Ʒ>4N��½u���A�=��l��	�� u�B�a���J���>�|�ߔ��A�yo�қK��bMt�8��GN��n��%>�0ҧ��u8^�Q�b�~��I�!��e�|(ј����'��䌰�ckfy���ĩd
��?Rv}��,q}KW?�@��)�B�5�>�$H��#_�G�PD��'�HJ|��5M~�I����z��&�
<S
8`��pY�[��p<��^�aDzTC�M�0;�*��`���{n��:�5���@O����k�j��D��ih��B�L(�ܓK�d)�`F�s��|�ƚ��&�O�E��EnL�g���V��ư��2�Q#�w %��9̛Tm�:#~߄pf��K�_"��94��bo�u@���ǝ氆��oOa^J+Q[O��6�����Oo��V�$S��:pc��7]sf��
1�"�k��]������@��+���t�����;_�4U�Y�}����A�~Yy��zʅ!׵���`��S#�D�z��0!�S`��!cKl�t��ب��]���OX# ��H�Ǐ����.�w!�/��QC���D6����> UЛ�4^i~�63�VU���$�޷����V_H���f�t��
#y���C�";5��]e�!��X�$rEѲ��F�����L��+���6	�T��
+��Gx2�:���%X�;�^���:~X����L[f��I�����=a��]�ظY��Þ��]Ƒ���p./��A�B����%7����JO~?����ɽ򛟘�K%�?��ޱ�`����EJ��&)s���qտV&z`f�:�� i��E��1}C{�y��b�7-�eO�M+yAD����PgDs��g:���-)Ԕ�O۹�ꡓ��e�<h��D��dڪ��4'������
��[\�4��6��.mYn�JE�1��)�%�l��{j�J���.�*R{�y��D�4�@�>q%w���7w�BQ6.ݼ��R崆�t�		1�%g��`�@=�{;�jn&3ik�S[Wb��}#u�"�/�X:�ܽ.TOe�E��xw����Yu�k�g�Ob>�Q��߄+g�ߝ�)� ��� �*;�7[ay�%�z�C�/���/�=��+��:���swŅ��2<����Hc�$�2�����<�(ȹ����4�,��D�U��gic h)�<N!%O��u}ۚ��J�TN=�����~f��ъ*��UB'�v;%?������ҝ�@e�5?��`x�c���c�g�����yd�[7��kF�O�[�&5����Ĝ�/�	�'�r��Fp��
�b+!I<����M���W�,J�yd^?��w- ��7:3�jyW�~�m��?�>7�Σ���|�{�D�Q
��bYr���q����"�'�����;a�"d�=�U��Cze*5ůΖ�(ۺ��@��0�dV�1�H��t��F��I��L��_�|�Q���Ҹ�xM������l��C�Y�
��ߜzB5�*.(i�u Y]�����G������g#;1�Q��u�.y�o�L3�O'��Tѥc��.��b����!�*��=�2�jy5,
�@Yʫ��m��^P���@CO�X@���H'�^�QX�[�dW�V��v݊���:�Z�v�$�/�ع7s�� �H͕Lfp�>���`>��XQ��*���\F�1�P�`��>
�p�Maq���_���9�$�r�Ē��ۡ�B��K�~¥R�����c��Y�p�}7�QB�	��2��Upֵߊ6U����۶����ڍv��c촷����X佊�d8����p`���Ȍu=q?��^zh�x	����1�C���I���]r���mo�e��qUf�%^�ʠ!��6�[~o"K� m�<B���-�<4�+4�<�j�Ew��-��(�i��}}�\�*����������
�G=?8Q±��e�MW���M� =m�U�3Kߜt�ڕ��o���۱�Ԕ��FL���9��^��� <�L��k���R��j����w��W�*��1��i���S)4���O��?"E��0z���?�U�Ql�Q�X�i�����f��Z�X	_��g	�1sX�m�1�o�:��kn��r�����K\�5x��՝r��������Ga�����mZ>r�:]��c�/��@f�Ƃ(��Tަ_�yyQwr^!��]��T>�"k�Y_��D�d�~	/�\P@��~�S�iJ�Ml(������bAoA��7�f< �+gS؇�Dc4 �� ��G���G����oزWGK~w���Hh�S��U�����k�<~l�r�?9�r5G�S3��9���f��N�!�G��49��4�-Iǥ�;����:���V�cN�F)�=�ť���ʾ~��X2�m�И��O��;�!�x̾��i@o.1�ǩfcC$OC�?����j?�$Y�~�1���8C�2���z������$��-!k���#�N0AT�zl��^�V�qj8�2�!�{btztWs
Q���Ji0D,����8V����7�iဣ.���R������~Ƥǌ�*��?�S�	�m�����?���Wշ�qG֓4=�[�؈����6�%E���.�m�.2��0���׷�ӛ�)|�h���ɹV4<����|t�x=̋�rI��qg`>SD��55��ޜ�h�oӘ��c"��J܉����o@ů��x~(�=4�&\��Ki�����Sl�X�].܂����]߲?�qY��@����GD��3]n1��O�9�Jl�����n�A�9m����r�/�[�P���;��u�G5����p6V�WDR!ң[\X"G;�P�S��p����d^T�ϐ��2��\�A���_U7"�3��ӛ��h�Ci:�=�m2��p��-�N�;����[E�L��Ґ�P��@Z�
,�dŃ݇�����E�,�,�<�'�Y_y����Qfrc|�����qz��{_�[��n�a���4�:W�+ �Q��3�}�����GX/�Ut[2��s�_�r�!�⥻IP���E٦�AUS���I!5�Bٙl�l�bz��P&�3��ݧW���j��ò������G%���~���X�*�a�LP�](�c2���a|8}+�y���5�Tr�q�uWe5�.���Mc�a���8z}"L����w�EWA~�Z9�c��2A�ݡԋ���M)=?��'��2Īw�.F]
�G�OC�@�5����V��#9>P�?D!�Nt�*r�>�i=9Ҙ�����1DF�����YJJ]�|Rd�H�4�u��8�o��U��e.���א����* �����Y�/J�F�{�MY=�I�'_�Kc�q�i(�Y��V�����;!$E�XɟC�b%���B�HC��#0��f̽[zm��.&�
�t�KS�(��F/��?]��q>��/f!&9�~P<��\�H ����-x�
8}�u'�n�����[�����4)੍{��a�o�O��X��{|���(�}Ba:Z��z�Gm���b)rem^�+�zrG\�t��.{�J����B�� {e@֧}G�� �T�p1��A_�3��KWIbzӸ�ʰ���}�>ң��25# ����&��Q���
�jvGS�Nu=���&Iϣ@[j�z=w�0��ҳ5B�%2���h��5*Z)A��y�i��M�������ܕ�"���5${�aN�U/j@B���z
f�?iUsH�b0B���B]Y��ꥶS.��m��<U�
[��U���7^gcz{���W.��|��h�I�w�$�g��.�a�TX}�d4<:��L8�}��.���}o��P������0*z�Ai�z��;��hژ�:��UG�z1K��2���\ΠQV]������=�L����{.4���������a����rl��3r�X�����¶(�M�p��뒾{�D1�؀��A�	��wa7�T���.�*�k�}*�o��rp5��	���b<�sb�i����µn�!b	��V�AU��sP���r�=���#�1*I�}f~��ɗZ��0N�S��_�9� ��=� *��i�"Xj@� .����i���%O�m�/�q�4g�_Ѫ�m��i?|7#-�g����Ec�hg�Wf\5%�+�G2�&��z���> kI�C����
X�K�8�;L���)I���n�)��j�-��Tu�GKIp�������/7��*ł���E��^r\K�t�ʁ.��n�Ì�n�n"-��ˑe���ꡐ\�h���Q�)�3�*i��V㢉�퇹0	M,ݖ��>�2���
S��[gt��E9e�խ�ʩ$���?�i�,4{��r8���X؟⯨�+�dÖF�T^��4�D!��i��|�ɑ2�=�%�Iٴ3*zjQ' $"H>I]�m��QT4�ͩ�$��%�|fH��;S�H1��wuD�
ĵ��|15VV�B�&c�m�*�m�lJLMܻaґs?��JOj%	e�6�CP� ��T��Y���X�~�E��I�Ȓ�gOB
[��cS��
l6H�y��f�!��I�ۓ�'o�R���dE���E�)-�7���|��\�H;ީ�5V`� $>�3-}4�*�<��f�e4[����O���w]8����I7�>�d�w�S��
��y�"]畖n��)�^$�
��f�tT���������C�V�y���~��K�T�]�p�24�=�'yG�g����E���� }m�"J�Y�x"�q Wd^���(����uL�E�ՙ^�gO��Ӷ���DD��AB8Y>cG�43�d{a�-o?MEץD�m�>��W�v�,��I�~�#�rG˺���V$��ޱ≑�	Z(�,�UqШSb���X'��;�5�AC�g�/��dZ�6�� �l1w�:���V�F�x�_w�UEI��� ;}���n9QI�=�Φt�
1�f#������z#߅J�qű�9Cv�+`�6�u�����ζ�Ե���^Vu@���v8��j!:)m\��j�'�!_��b^�m�R{�h�-G��ƎvO"��v<Dz�4�`�$W��v$���䒓����7��k���IQx���"o_,96Z=<�j���%�-�� �n&����ڞ���7[_bt�4~�O2���[!��5ɳ�=���$QdZ��@3!>j��Q��/�6�0�<��ܪ�!�ǈ�c����C�83m��1>���M�«u@�d�<�G1Lo��#Y��ӑ�����@��t��t gO>��V7��
�ZIj�6���75a�~:��	Yb���[�5��U����o@�.ĭ1�V�|τ�pLj� љ�o�q�ՖYDG*����y9F8i}M�~uOP�q��#�� ˶R��r��,��fe+i	�I��|D���t���H Pn��</�q��Фgi�n� 1��q��ў�R(ɲ��km0�V��yJ�pJ<�{r{���R���QX.�o�����m�R�ҥ1���h��g�8�Ĕǹ��t���8�A)r�3�
҉�uU�"�1�;yP@L<��2B��\�\<��v|>��
����ŵV5�G���@�_jc�҆���֍V���Pc���ξ���Q�&[N�⛩�j���X�O%�>m�E1�k�!�0�Ʈ���3ۓ{��M�@E&�ꛬi�Z�Ck1g�H�;��=��w� �/h�V��Hs>&�M�樎(}SF|%����j�fy3�c�F(�/Xw�С�7E^�@�rҌ;�G8��$����~Ik�Z>�a��s~��'N�H�f$��;�
&���gx�OY\L�L֟�{�ďm��P���>��G�?�C�5��d0�A�V��\i?�X�
��Q~��	�M���fcf��5�d��px���ŋ6�4��ÿ��@u��׾Oh-o�JxM~�G���R�O�$=3�f�U��'0�#�8a�sU�����X5]\��>�gr�s1�O��晸KQ�{5����7�Q����%:�9AF�lPC��k��SI0^���?Ca�\��͉?�0Ս��u��>}T���w/�1۽�u�*�1�P�"���y����m�ģL��e`��%g��T�^Y�,��Fҽ���*�x�Χʢ_���/Mz��K[��3J�J��a�ȭ�U���{�*A��^�o�u48܀��w-���W1����-���<��"����z�6�#��rW�����a�o|�)��S����<Wxq�^q�dy��|)l{UV�{ry��[���'
��3�@�G�AARN��܅�􃹮�v[nѣoKl	[����_A�3�U�;�{[���Rpc��+��:T�,��L$��*w�M�D�6EXlɶđ�S��P�9d��hgC�/���`΢؃���0H��MC������)3��^k'�KL�Z�:yj��/�oߌC}�^ 1��m鰄��;J�`�?�����-qh����.ԎK�����,}�w#x3���a(�ꥴ�g�ޭ����x�o����c]�Ӕ��帪|M�`/B'�8I�:���!A%ꌏ�
��]�����c��<�a��s٘�FP�������}	�C[��1�A���7�f��E�e���i�v�ıvWM�v'uל�1�0�՗��[18(B�� ��Y���s�o+�I��1�F�**�p�9B�h���}3Rc
�J6}�.g���'k�ST1�E�%����s�魧o��}ngJ!Э=I�V3��K�	ew6�,K�3Z�xF��}�\��e�k6<&B\�&��7�w<���t�`�Ue26 � �O�a�}�̊�pg�b��Oi�;�v������uxK�us�;do�G���1�3u�������7�KNM�͕�r�w�d|I�����C��N�w1��]��8�hڷ��-��@�_.T���H��HS��b�u_^�8�����KEen���,�?|���f�`�@~6ݘOxn���Vy�מ;_q���9�0�n5BNq'�<�8������c{���3�޸��3=K/�"3��e�t�M?�2�Ò���g3�9Ǳl�ґ��ɳ�Z�N��0L^t]s�H�;��a/ֈ���S.(Yz��0.'�Y�!Q�^�C^�r�jqX�u�	�lݾ8(޵�b� �H�1j��o[���,�-s�ڍ����kߙU��$V��Ft�=c3�y߆�X	Mb���M���4\�^�����Q�ܸO&�l}��a��=N6��[[�DS;��j;��/Lٴ�M�򳬢������@�����G�[H����gċ
I��lm�?1ռ��6�G�#�	������c�V�ۋM�h�O!�H(_!g�E��6� ��c�0,I��q���j�;�2N��D8�4dZ1�G;] ��8ɢKc
�R��*���fs����X]��C�8���:n�����$��PA:Y�m*���{�ڦ���v���1���;�b��NS�#v�n������gSHf��<
h��
����<��*%���Caf$�����$��<
��q�4���ZVq$K��Զ�.�Ry$m���9����s<~�h�E+�z��1o:�q��$i�r�	9�5�Əvd�G��"�}��>b��'X$�yۨi��,�/ǁn�P��M��O�Ƚ\����h��V�/zS|Ds�����Y���AʸݽN=��\ūy�\G6֞�F�
_s��Lc�gq��0�%�M￥��5bP�t��GDR.
f�FC��³��fPp�^(FG�HΓ@���U�O��Jlo��j̌,1㌥����1Z�j\}��Y�^%�����Ρ�Щ)}d �8)o{E���%���� v�R�6c��c��}��U�,f���6��^������ق�@ΫVe�i���@=�����n��Fe3i���M�T�Y2�U*�(�̉
�Iy	<-:���b�7�Dd�BU�!�~&aޅ���9�pi�+{�V � FZ����7�]QG�9 r��ڧ)�MA����RMld��N�'�P�8�y�,S�����Ω��V tibd4�C؟�'�zֻx��j�m$�C3��[���n�W4��S���F0�%��^>� ��Ԑ��:Њ��ud��䨍��pW�
�ۤۄ��~T{0d�V6�@�W�/��泶S��5�9�Hq<�!.e���P^1�$@�/��<�*#�V���l�CH7��G�y�=�ݳ��W�+�\��ޜ��k��2��A*�|������0�7�û��p�D)�*h����5�T��I&98�܈/� u��Q����Ԩ�Z� �F#�"pɺ��3����O'��h6Ea���Pk{�rpF��[oT2v�A��(�ٽ�w�G��TҨ�9�����j�mkM�c�\�K��P �Lmʲ�g�\J�}��C�ȓ��~ہ�m��� e�h�_��w�{�����=�W�h+��Z�+���1&[l'$�>Z�}Ux��oEtrI�󕷏��r�f	��Fd[ �L�u��5��e�d`�t�xq>��n�)v�K�#4�����B ��D��f5�ylxI���v��H�sp���!i��x*S��&W0��n��}�iM�q0�9���O��E�� �V��6�1v���85<7e2{p�c�g�^���[�=��վ��4�H@��T@�m�n�)������'|�D2¸(���aOK�^:�������=p�;ud�rg�~������r���ș�l����M�~���㨮vZ����	
"�:4�:O����ݚ������V!�h~p�S-m�v��P��9 $ S�p^n�X b��۝hK:�:�{9Ļ��(~��*객���Њ���B�H��LT�bi�l�����Lg�ҁQ��T�O	!x&\"�;Ҝ�b�\�g�Y�'����/�,,��x�P�+%+�N���Q�GS2]_�t�������S䬺 ٘v+��(�%�;�	@�q����I�����I����s�����C�mm"��pm��MJ�������u]��i��c �gB�˭@	���\���9�6DQ#l����x��!-�������y�R8F
R��Ӷ0��fWIG���O��7�D��8x���-C� ���-e3�^��D�9����+�aꚖ�$y�[v=��>I��,����G�-����Ɓ	R����O��Q��lw��}P��~5#H�*<y^|6nK��gK�}7�������
T���T��ގ��)j��(��7��gi�2s|��3�����آ:׫}h��E��]yGV�����ģ�ҎR6M�:j��^��=�b�W�gxv�L0e��b@�x�o��S�}S��E�����j[D���r�^�2�ȳ�=H���Z\�=a4X-��p"�(�Ѯ&T�~��s܂��B�56)a�z��J�YY��Q��W��yb���_�T��s����F������L�͖��5�a�[�H�<�Ū�x/(we��������2��iQ�k?�A�R��	%���}�Tfٹ�pb����bH~?zR8G��W��ri��3�(�L�W���-� ��	�4�zqߩq�4ѐ/��bK��[l<a&:珋?X�vQ'�J�I��������f��q-X1����yU�,��P��.��]'ͳi�NT�Bٍ��H1�"���
��KHB��<�˔$�E����I8(���u�2����,w��)�KY�q�쇡�l��r�T�^������ka�S-�\ݣ��� �r.rv��
^W� ����lXq2�f�{�R���	vFZ�H;X���`���?���dQr-�Ks�5{<��pQ�D�/�C;YJ]�Ky��/�ݭ�
�T���y��2U��3�Wd�	A٭����j�A�.xF������� �B΅з.oR�T�T����]\�![�;ˑb�D+f�,��]�۱��׼����4��J�5�=�t��-���Ăn-�(P�x�x{|�E�'���&b���?i�R5,�~��IΌ���g�u���N@�\�8Ml���,�����#��.�����@ذ��}�&�� 3jsϐ��@��p\?e{q�q�k�+WP\�����)�K.���v5����௝ɰJY���~��؄��#���G|a�i{f�Nߔ7�t[��nC�w��0G���b�����G�C�%��S�sN�>J��"~��-{��ʅ|����@�Ml���SB�١�'�C�R����+3$��� oC�xXy��
����Ù�Tj}�]��q �]/���`�@2����4�	'&�����`�xj��
�z��Vu�5�9t��[i��y¥�P����@c1*Vӊ�CT�O����$������q�I�����)	���^���D'K���Ml���* ���R@�s:���˳WJ�,�C�\�e��ޭ2���hܙ�:4D��c���qt��u��4O��G��n9�a�~��Mi�Eٷp�_=�C�=�]4�A�Cl'��z1�bN�H�z`����]��~ӗ������	>��P4��Mg���D���{�Eu�s��*���q��\2��1�zkK�.5�::�Hoч���N1E͜���/H	:*�5qs��@�	��y��(~zp�ꤩC�E�:�^K�o�qٳ �Th�!����o�56{32w5�#�oS��@k��e���ؕ�غ�w��F͉]����#��g����l�H�M&�a��������,0 ��MΓ�v���*؎��R��*3���v��;������NK�����*&H@�H� ����������/Y���jǩH`�.v��z�t��\v��9�7Vx+�{���I�=p�����\�n�!#�>>h�;@H�H.!�oa�W�RP*�e�mj..�^fV܈WOn]R� f���.z�')4]�B��n�������ݓ,�t�K�s)h���wx0\�]V�c}�H��{x���A�5�q��x<qN�u��c·Z!*W[	��m�9���q��䂱��f� E�Ů�n|4%�[�APV@6�jUs����(�5b-��8ՆÄ��Z�@iU��ޏ���QsC���Uqn�����DF�5+�"a�G��'�zhؿ�u1�@� �p�xgf�H\�LBK��}4�zM��~��'�B��L� ��n�����e�eR]��\�#}r"Ck�U�AȌ'=\�޵�񳦏ᆣzs�φa��_ CF��d��	l� Y5�~\!�%�� ���Paĳ���c�,'c� ���k��A"��&��mG3 �� �d>���#Ȇ8��/S�"��q;������i٥��?�h��y�\V��88A�e29�#[\:���O�϶y�N�nbr���R�hM ���z(@� $/Ӊ˫0�wi�.� �&�/��[F�"ygj'#&�Jb�������$)Y�b)��[�Y�m����H�͆���y�ilV���������.�<�H*�qܢ�v ��\���ц�M��4�8\�4�����H�l�s�o���^�~�x��ekvT�#��'���`�k���%z�tD�yo���d!��̕��ˌ5'���^����g��TR��P��ůCd��̥��X5J
>,o]�4	�b�{#o�Υ�Ś���7�/_��$���^ݟ\+H�	kC ��}F+]�_���Z�oov��ic9Փk�9�a�����ֳ�.຦�͖Y&��MnCi��^��C
�@arn�F�\�F��?�����)!�~JX�Nj��Y�%-ul}�m��}�3��F�d��LR�u�lҰ�
G���nMD�J�
2���[�/�iv�#J�>m
2����f!�gP:q%��6�QO�̂<�q��5Vv*s�p5�s"���kє'����'���#�Z�����W��?�EX�)��G�-���6*x�~�;�:3S�GP8L�)?� ��B�����ѩ��+a&�,�9[l�qC9���
F��9� ���FqţB�g��>�D�~����_Z�6R���N���|���#|����?�]�Ȟ��U�D��0AL�"���ks ���q#&�{׼�TC�z;/&t�x�M�)ԻP|1��3*�R�_�);o[����9d�&~�� �d��rE�1�)�hG;w��l�Ov�
������WT=�lu�1�0���"�O��}�$����ΗQx����M�~�M�⑨�M4����7�h�'���X�UR�잗���I9��P������x��s���K�]��X���7��k�׫�b����vc�e��,�Z,������I��G��2ĉ}�*X�Y�	�璃����愈0TX\Z A����(��4��
�]�/	�+ U,�:Q!��ld�/�|�j[<���-jO"Lȁ&g`�G�����J#��9�Q0��!G�s��pE��L�T�_V�8.�>�	3�)�f]�S��"^�!�f�w����I��%F�%-����l�] 5�܇�v�rg��9);�nM{r����[/Ek\8��ص�d5� �\&Ύ��� 1Xc2����Z��*2
�~�qj:h��׳�2�k��[��g�F�� ���w�V$��yŴ���!_z��%���$�X����vZ�aZwqx�=J��(NE��_�'����e�Ȩ�f�H�Fq*=��L�QoQ��sP�!�DuH��
!��*%�d�l�^#!��R�����xZXw�oG���%����t�T_�A͹g����sH�[��V�@�5�	.r�DQ$l�����ɢ�B!�ˤ�婔u�^~���(�s��n��O�R�F�~5E�G�M���/��7�B�ى�&J���f���Iَ��	�a'��RZ
��7�E��?<߰��'P����q�}��[�(lս�Њ8a"��Hg��QAo����6؆�7N�8a��߯\1���}m��b4��b������!�O�#�渌�`jMeDd�=�m����[Ϻ��fw���c�oA"�ve2�������gi��Qz��k�qǐ��C�ID��LW�Ik��ifd����:N�H(C�y�����F��F_�FK��.�N��)R�#t��#X�i9�t4U�4rP���[{�a�AY�c���@�5��ta0�4���;8����W�"�8n�@}@嗲����yJ�6A�ۃP�7�K�nU�h���qAeO^�^D�Ț���ۋ�1:Z)#̉#ix.7z
2�h�S"p$G����Y���yq��7	nX���<�l��)��RhD�1���邘\��G��SvE�����@����خ'�V�t.�<��8A��^��(G�#6�q��~ȅL_����X�w�G��|AǪ0�N	��%����`���2����s�R�V"ܭ��'��'�']z'�t-�-w���%�� ��#�T�= 
t�h�Y���/#������V��/���c���2���/�c���j���WH��`\'�E7{^؊�D#!�mt��z0$����{��.�~�O��^��Us\��[��$2{��g�I�nnX�䂏�5�]�A�lP��զ�&1�;�
M��O�j���{*�$6[h�Fᯥ�x.�ok1+��G/*QR��zӦ=jU�i���x���|!��A"�I	w�Z	�tLn����i���̌R����f�������#+8��]ֺW���SEqڌ�^���v~�nI�A ֙*D��Y|�r7н�H��s��K�zro	#拲���
T�m
u�%���*�*�O��޳��a�}h�a����9b՛�m��J�:�ڤW�n#�*[ض�C�y����+��
��+�XlRܑtޭ\�wT��D&�������K4z�k��!�&����9;�U�?�U{K�@�ۄfhx�HP�X��f���P��J7z�3��qH��8f�W�Ư�>�^�q^��H����J�V�`�l�$��A#��w��|p!�3�"E�sv�;�>���}��oU�x��!�*��	-���}�u��<�F�;R�Dh����QR���K{.[�6���a=��;��j��H��	j����/�����LS���#��M,-��#��|�ӈ3��<*�B�n�2W�����
��	nJ���;���v��'Cw�.��ݴ"��w[��P�R_ �;^T��2,��NI� +¬����94PAt�fD���&VX�vn���ț�j�>L�"U3��7�D�~M:g�����$��������0�����pM�+3|p ݅t�l���2{WIŘ���`�8�z��5�'��ނB]v}��5x��E��=�5m
M�^y�2ۦ��C�仑��dY`D�
>?o�;h?�\z��^�Ѱ|g�.G����'3��}�B�8�8s��zSۖ �sLUI���7���M2Xam��%�E�X�=��V�������d�_��p2��p}�gCZ�]�dSmV�����Kӌ�D&�w�0W�u2�����:��Z��H_z��&^-�L�f��y����X�D@��n���F�����\��)�p���$ލt�:�����/�>��kΩ���=��on�p�/��I���<@���xN�2Q�ejΝ[�>N�I��xA�Q�KK?�*��Pv P�i�ԧg�E[0!��U�`![�Y�Aҥ_�9��(��=O&�ļK�݊K�? ��!s�?�d�X����>�	X�5o��d�!Ǥ���U��V;\�Xl��@��*Ȋ:���V��l�����I���L���oT���E�H�Ow@('�WҸ�6��h=�������S��Z
 �q���jzQZ�.)���<���݌va8���X�>`g��0AstŤ�z��يdT75�g!�g��U�)a�wL���6���7��KȔ�,Z.�{�xe}c���W8�^!�0�z��BнS�5$�
�CB�����7�qU�t���J�rV��Ld,��~�R$+���˨��!R.�0��齣Ug�<�Ys����рM��:ŵ����6�nP{��/�qq�ώ�.�_y���B��^9qh��������9H^/g*I
&iO�\���>�K7�^�C��7�;�;�Aza�@���,�*�O��^TF���YB�A/`&� [#h°�ٖ1���b�6m�减vBvrDS�Q�-�;�8d�\��s���vv'�o-������¯(��U�E��ې�Q�_�����>����mh�IegxO�a�<�~�R���.o��}�g�z<���7�%ki��Ʉ�8����R��=�%�_��I����ZrCw���$y^���BTyA�ɒ��?A���M�t���@2�c�G�$u">�\D֑\EU/�9_Nb�+,o�5�_aEz�;c;�ݤ�4Wc�PA�<X���\;4
mm�k�~�	�>x�t������P��x`���B���Cp[3����g���̸����sac[��
I�*���)�������QA���;{AJ��=�6�`��5����>
бs��%��P��e2�pn��tCo���T�"Č�E�
PE�H},QY��w�'<�`�8�/w��O���E���E�}��(9�a|Fݿ�a��$�?4�\��=�8�a�+w�z�ƺ=��a  ��d����6f�=R��0˗����Ŭ���^�7��)�/%���(o�\l	{Bvv��������H�����\v�;���i��ˮ�k%��rl&��	<})��1$��Jσ3�V�N�����"[�Z[��+�P�Y���2��9_\����Ubथp7�邋�,�V߲BKQ[�kɱ������̾�k�4T b�����{q���@��5ǻ`�i�}r�J;2��w�}̯�٥��{Zw"����2�H=l7$ g�<hV�a�����I�\Cx�eJ�s��?�����wqBDz�c�b?�{�	Z̼�u5F��v|��M�kF=x~�c�kR��*�����q:���n��{z{Z����E��s����"m���İL"Ĉ��#'+!�uϨ���T�a�+.Q�3��2�r�(�Ǟ>�3:��^�$B2��T9L�R�*TF��:�8`yKSթ;�ʊ9X���/��ZS��k��*\�jﮄȫ񠪈n;���D���v�u݋��2z'��+�G{� E��]�?L­i�4���[�f�Q&Cвx��3�37f�C�Q��u�0�$֧�$	t"��(�C����~��o��Y$,)����U,M��5<FI�PB�y����R��[-T �V6�ov7
����?pfA�|ڛ�h7���E@��@w���R�HZ������$YW�ǪJ�AE#(�ik�/��w� v�����U1�2��: ��_ϞJ���*�A��m�,(U)�NLyj/���S��m}c� �*̄D���d�Vߓ���N@�`�-�ec�nD�L�D�ǻ�Ť@B���$�p��XmE�p�m�觾��yA���	[A/�D��Y/͘�M�,0�OFe�Ș��|�a7Pf�aR��{\�:�Z�C����� ��X�M��z<.�؆V�8w�:��oX0�0P ��+���g��h�i���|���~���(��!��Y�"·]e�;���.�v?Q8��n�Mi#�&�&�]���
��J�䫘g9��Ġ���ݽb�f�+������S�o��o�ruЧ�C�x�p)���ݩ'�5� �	}ej���/��r>�=A�K�� C���MT�L`�7C��m�����?P\y�b'�3�\�!�,c~ D��������~�5}�&�V6�����cļA��5�,?l�^(M����
�44��T#��ȱ�D�?���Ԙ��r[�OtE��`��k$�[{��cIP���(?{��P�K|:E�=`_��w��Mg;Q�^fZ��S�� Ā�=�rOn)���)oO'�G꠸�8Rٔ�0@�;2\�ׯ��w�K�i?iXd�  ��}z��6��d������dZ�/��?a\W����d��3�d�+:$Y�S�~��"�;��걀%Db��p �,�W����@ ���OB7��.���+��Ւf��n?����F]�1l��������&%-P�2'�Em�xZ�|B�S2��S��.`謝��D)ZetC[�L|%D��}qv;`U�[j�6\��4�����A����G 1�R�c�RF�Z��;���<��E�� t|�iƾ�'���ᑖt4��*Q��a#�M*lM)����GO�|�J��#
X	BA��}s�T������M�	��D���~��¯�|O_A�Xڏ�g�샢)���qO祶�ӧ3��`�̸ȉ�m�x�Gs.��0�C��d w��$2G�0��L�Y�����.��Z�$��"7�Ugl�pDy�Ӑ���9�Lh��Y�����
w8��{��+�׮ݵ��k������kb�;�m��G�zH��8i}����h��lE��f.U��[?^.��r{���}o�5M�{�D����������:T��ejn�6!�qZ�d�,��P�d�&o�3;���}�>�$��r��8F��F$��V�	��t�ށ<Gί%��b ^�/�{i�\�X���+�$;$V�I����Պ�~�ˊ<z��`؋`2�кq����ƁW��e��p�.�9_��Uр��Ac��k�a�����G���b�S��Z��G�d���b����Y�W�'�0T<:d�L��g�Nwx�楕%�/��zh����)
9s�[�� >yQz�GK:�`��Z����£?��0]板w�ݝI;"�0�j�x#A%ɴ��i�ĸ��T�3|t%J)�T��J�!��P�#�$��Kᐓz�#�j7�@Џh7��'����`�Ȣ�$��Г�yT�ٕv>|y]ΝL��T���M�S�E�UQ�U��/�Ԫ�T֎� H��Y9�A �����d`A��Jx,�9aL��N��hQQ9g�Y@Ƅ�ܰ:[�z;����;,(�����Մy>�������z�he�e�j��5T仵*��U �ɩ.��?:v+��˪ߢ�Ƨ��^�))@�r.`���,o
��)|�r��(nnL��@L����c�r��/^�ܧm?`(V�n��%��i��jS o.�n�{�=���D�AH������CQ�L��_�#$��ֻ�����Ӛr",��.�F�#�w�5�������RtL���Q��ab�䎫��7����k�)��^��8��@H�oA���v1�CRR���\��c���{�,ը������Gp�����sd����朙l_B�0#.9C��q�DY���mڕ�hb�K��㦺����\
�YT)����`e8acA#H8~��,�^uK4Ci���u�}�t���7#;��;����(����-�WA�Y�;�hZ�c�k�8t�C�Di�5!�#\��+��x������{�H�pYk"���^lb/Kph�`D�zآ��&�{3�<=P�^h��o����%ᐌ��g��x5���gb9I�X��
�O1��ќ�D'�i�w ē�6��-_�~�Eã���h�n:#`�x�%툏˼��x>�w�нukՀ� �I��ۗv	&�61b�����.�������f�Y9f&�A �S~�� �Q(KD��e7ĲO@d�ҟ��r~�`��s�y�1�hx~L�Gx�>�S?^b���L%��{�����i�������P���H<퍨u����PW%6y�i��L��k�O�q�����^��\=��cen�@�{W��Q�C��Uj��� �(;��R!a�͉$��߻�4�fT|��\��Z(���q��lx��s�T����_��Q��ؾ4�{�P�	w�r�@���'ͺWD��W��c	����R����N�i[��,g|�}F��G�GD��[YaqG�<�\t�����o�W��ٯB4���"5�O��E��i��wqc/4eg��X�eߺ%�8�S[<P^Is2���k/nD`'�<bDΡZ�x>�<d_C����u'[��){=����B�>�?`D���0������.��Nů2P����ig"a���Q�tQ�	���)z��`������˺�ДkOT���V�IP*�f��1��#`���b�"Y� -;ʙ���Cu�j�U�w���H3��b�n	c����Ss	2bA9z�F��c�e`r�=1�;WJ��Fl�Yk$��To�/�������Q� ~���RC}���V�r<�q��Ca^L ��ąN�N�[3YA�їpa����o�;�B���������P�v�;��\1��^\��(�/�!�#�T��*T�b"}��u�d���]FjY��V�]aGsO%�wiB��E&���$MV;�z�>=����z�T<�ON�Z������ ��/���z ��:)�>ØʜN��e��+���܇O�����!�y���Y�R�gL/3��n���˧LT%כ0������}$E�Z2�z�,�Q�I1��/_�@������ް�R/���CC�qcE�04�7B��,<+�d��_&�딗��v����q�K$�y�	�>]�͟��]��P��^9ɭ���9����Rk���wj�H.�S&�
���N?�n��������'�,��Ж"�G���9'`9�������: B�R�$5l8���]&��� ���S�Q�ӣߜoo��Mo��u#��y ��8s��ɢ�1�#_�X}P�Xr.��:�4EA!_����#���o�]��m�] �;p�zڑ��7W���{����dq���aXi���/�f��N�@���~ߗ��� s�V��`�۴Wp���w�{��L��H�)F�#�^Gg��,[.9�9OV�r�E�^e� �����a�٭	K4g�d����u�*Uu�n�E/�¨��j-��5�L����_��ji�^������v��Kȉ�4��
7��?7!-_	�*��%��cL����Z����3�8n;�HY�t-�)�p�{Ѝ�7BJ�v=��7't��-�� -�U�"4���Czt����³F�o�T��q�/����[##��c��W�UIo����4���("a��Ԋ�vtSm,J��5��9_$P� h����B����q >A)���z��3�]����̩��6_����y���ـg�zQ��ջ��yW�(�G	���0w�Z�,�6^�:z�%W8b�E0��1����f������Ď��Jc�#�h^%�_7���b7����7XjU,{|D5cs��ZV�Ă@�to����T�4���+0�:P��R�rd����c;�Ljg��Cs�=H��v���Ҡ��#&�j��L�y��u#�Ej8u��Ͼ(����rץ|CS=��e'�OV.t�Q!��X�Y�[
�h�P���4�o��g�D�)
d�f�R�p��.�TO����(�o##�2�F��X����V���M`h�{�q��h� ���ћ�7��e�-z�,���9��wJ82�u��X#I�p�/���$L�����K�N��I��
׾�W�&QަOʵ��6;��N"��yoH&P(e��?o�K?.	�N�_q��ֽ��}`�7��)�&9.�������ϴǵh���w��s��QB��\��'��g��0Z�Ҭ����ψ��"-��q�I�-�C2D�|�E�y2[@0]�S�o���+�;C�L3$���M��_(�yDxHT�"�Y�j�H�?7���Fm6;�E3Dg# x�^M�5U�i�x����������;�(�}z���'��
�J]����?���%v��~��V ���&��[��/'�P��� ��4�dj�%�,lbAy�;B���;�&�}ė��g���Uߣ9�u�Z�p*�K�Ћ�Ev�U#3����_EN�@m�uU~/m���s�k�m1p��|"��d�A�`�+I�3Lu�"��Qd�
�����-��G[d.���Q�#�9�֖��
��W��Wgn͍�7T��/�>���:zc�Y7.�}�P��Kø:��7����ⱐ�9�Ma[+����k�J�����"P[V(ry�ݸ,�U�Bz�܉����ư����3�7�ךU�I��gq�Ә-2KD�e�b��ou\�vM�������m���t��� ۉʠ%(�	$q���x��~�C>9+�T�9mra�+�p������B<~N�ȭ�&�]����4 �Ţ� $B�EԐ��D{�R�5��l�pk�=�7��8rGn3�j�5�A�W�k+���Ǯ���c0t�z��5Ζ�h��|a�W�#�+�'�\�We��za�<�-���׹�}�rW�1켻���o��loQ�#A�&�v��.ߊ_�$��_%����l�Km��0�/�2W�.݇L
SY\�^d���MlRtt���)ax������l�k�jB3�>c�CAK��<�}�s�A
$%zؑ�T���C4z��:p�,��MҐ��P�M�.K�L=ؙs/���c��L� ��1ޖ_AV��MUL��nwd�,`��^����y����R0�C1��N��Ay�!!X��%�1�����u1F`��Nq��?)�5�eUzo.��=W��0��|�}t��X�b�EC[	�����p1:��V��>U�7-v���cQ�U4^��&=K��I?l����`�Y
@^3�A3Z,��͛��f��7�����46��/��'1ih&鵲Q�ظ*�-��+�i���f֘ԫ�c��"�o�� ��j�#�v�+=>L��t
Ѣ�!9x�߆ԍu������1lC(���u�{aO�h��6�$��d6D&�кz���]��go��� G��PzZ��+�;�F�v��|U 0.d'a� �
�\#,��zQ�}�H���m��Ήh��Ȑ����G��l;@H�$�>O��T�����LH���*ͨ�Kk����=�G;	��CW;�Z*d(�j���'���5*)�co� ��i �Ĉ�3z�um�[|��Mo:@ �^�6�y#9J쳇J�p�:�q����B��#��4��؜d�����&��G�5^Ù�;x�� �� V�հ��_=�� 8K��Ou��zA3�eݺ��!��������A�˰�����	'���u��c��}z蟢����E�$���|�缓Eѻ����w�Ή�h�E>b�O�|E<�yIq: ؞R /�T$oS_�xH��J�e(
���.Q0.I"�>)��Va�m����!dʊ���`9�c)(�����w>(߷�N=��tk��IT?ӡ��T%�20��B���v��s,��׮���X��6�M��[$]�q�١!�p�'��6q����U�q���Tk��V"Wa1�)��+?T�"4��7U��B�ݏV�B�b�l���hI�_[��P���ĭq�O ��ꃊ6�窧�,N��M�������袍�eJ��8 �J���-`Ta���-�O:�UN8@1|�	5��1lC��qc�3>����<-��~Ėxc�����w��o@����3�3��2��y���î:ɸt
�Z����~>�Aut�xR'�[���e� ��9���2���H�����=����i=I�h�e��0L�3R��D���,���O�A�H��%Ɩ`2]5c켗� ��Uz�j��i�m����vGz�~�
Vmx����=������uEC܈m�	��}�2����n_�O��q ��y軘�b�/?��s~���J&��,S��-M
��V>kdJ���ւ�=��+fp�ٶH����6�X����a�Vn���� ���15��"r-B��z�:�ξ��0��|�&j�{j~N>*M�P s���?jf\��O�E� ���7�P�����c�A���S�����R���M�Q�e�l������6b㒑ZV�.}��	㿱YE����rܱ���
�WI���&$��lN+=)M��f�o 6����
��N4���/"rS�������j��ş&����iU�7�C<��B���b��=�La�b�$Ϥ��X�2K;������a����2�GO���r�W���cB[qe��~��d���%���k%JŅcAF��b�6�`{{��:�l��d�>mZ��H�'���<��P��|��2�B���Z��/p�%���saW��7��g]�T�˘�~:�P��3k>,d��'��ǟdܦ�8'��Z�c�DQh4ck�-kBφ,E�S0�]i�_s3���-�{�p\ꇀ��8��ero]����$��o [��ِ
�1<�Րn���nȕ��N���+`��]Ò��*�#
�����*|y+dGr8XtH�Gr�tN��i�Yt���\�҇�p3�{Ο�0-8�����-!�kx�W���sG�4�XCk�Z��t����Y�E��'�Zaa�dYP@�m{���[4��V	]��|u��G�'%�sLtq�n:��!Hb�{J:�sc;�T;-3z$��B?Ũ�7Y	�{)޿b���~����(s�)s�9�>Wh0��^�5y]>+���@3��Ό��s�a3�}e�߽���a\Ͳ��=�����4��u�>�R�H/�����f��>�t�l�� ����B4-�{/�83�2�o(��m�lZ����K����d��	@�H�q�&t��ا�w����ܩ�������PΏ�����z���:��l!Ҏ����pe��T�^���Eu�# ��	�b�k�N΢ϐ�l��z	"�ء��P9��D����Q��=7�8cE�k�Y�Ǜ<|���N&�jDfxlql�^!m𧸹ƙ��+d����oGŚ�&�
�A�ez��*N�©�6K�J��y9"��#s��e��3���!%ɶч�`�܈f� @�鈗�G�ѷh �Z������Li@"m�<(}q}�-!>!0D7�DD��Du����4*��ї�Q)���������#���s��<D�2k"�OHǧb$���"�ԜI�-�F��@�ޡ2�����d=�G �p�W��_dgOgr�U����ӷ8�v���^O0���E.���T����X����/���$��6��5�3����^�q�;��Ps	�# Mu��;c�vR�^?�:�]�L��TI�p����cuj%6����,9�'E���(��j��ߝK�?�^��U�l� ��T�A�}�2���9�� P*���P��|���	�S���D�3�#c6Gk5]Yǘ�tN���Su��xbT�	I9O��9���I���c����V�������@��`fMI-��$�>[	����Sa_�Ss� ���#�����d]:w
g�������O�zкK{	 md->Ih�F BO��l�@ ���'���2(?�0u�$��c�x=c?�h��c�h�h0����v9���9�)v|�'% L�N��d��!+C�j�/6�VN�i��+p���t��u �S��o_�����P%�<q�g0��%�f��ۚU�TC�D��X�m����<�x��4���GY(n�W�A��-�q�?n�٧[ѵ��GԱȁ���u�$�9/�6Ȗ>!�Z⃅������
��oô�z+/�4�XFH�zjn)	��o�s������	���$q<�zu}���eh]v���g�Kg�ө�r�S��F�ǮNl�`5)6(r�!,�:�$n�0���=kPX�T�mC�LN�$�9L��	:�����}���,�\�C�Z�P1��:d����� X�T.\͈R��ʣWF�7���!;���j���]�<�����)7M��&6V(v:=��49Q�G����l�n*�F��l��Mէ��a��7�.�� q%��'�J��p���lf� �fLV�x�K�6~�bp�@��T��r��1�x���������"w�W*iM@JC��eT@���6o�ay�8�U�(�ҟ������|䞴�L^��6�������>t�*T4�/E?FO{5x9�sNWqp��*1Z�H�i��>]��6��H��1D��-%��O���;E�Q���1Ġ_JRLv )���^����"b�0j��p�w�[I���s+�L�}��"���c���m�n?w�Q@�A\��������~X���3��e�0�Uō�89$�\8)��T����2R��s��*f��!l^e�z`��cZ˽r�������NF���γԩ��K��St>�#/�V�.�K��6?a���v���ס�ϼ^@o�&�{H��g!-\���O��S���?�ށ�c�;�Z:Vǃ���.���H��ْ<}�����!�o_��a=��]�Ԅx4-��k���41lEr���Y���a�N����A�D�^�D�v!�U��O���v�Y�%�\�L�#�hz�:f�h�W$�p"^��Ska3�X$ǔ�������a��h���?�C�6����*��`�(QvN
�����@L��;��jT �<�7{��&R�CB3�@�C�4F��^LU{�$#t���(�\{2]W���7!7#�M��pۖ��j/�F'˜��>�	��j�A�:�U]�3pq5)����D�n_%[�G��)]Ə��jTX8Գ�'����.�D�h.	T�����P��*�t����O����MfQ�������=�re�m�"'L?�1�"0�k(	�`8�ZwCn���$s�iV�H~g�>yk1Ӷ�} RJ�z���G�Q���M!y���������\ 2��r��O�����w)��ɂ��o��Q@��z;
"�>0��!��=�)�K��5��B��xzZJ�f�TȋhC�y��u
��,�o����+-cc��
J�&����ۢ-lF�P�L-����ĀiLT�f'х�q����0~�L@?xn��8˼t��S���A<�k���c��McԨ�E�G'��4��-��|JR��-��!�Vz�� I<������h�Z@��z0$�Q�7�[d�k����&���\DTu����@aUU�$��H�%L4-L|�?/[�ź[�k,;��mH2r	�Q�m��R�:��0���!W��'UWuc�A����N��lwSZD�b�q)�L�K�ZPU��_�`�dy�d�W4`�����f�	�"��=����c�̬{}Gaԣ�!�w��W��3���"��y��C[F_��X�O"��+�I��n��ixJ��6���Q�t�w�[�{}z�LD �׍6�BUa|�E�J� ���䠛�u�� \��߭�e��U���#�_:�{�K�̋-�Am74U�ve����%�nAs��\���3��:����r5l�ڭ�M�Li"��|}����u��394U��9+����z�诏���bJ�9��o��2�T�M�?`�p�_�d����ƅ��e��%ȕ�}��j�
���-�%��xI�5������,��{䤧�G1�ֻj>����"|�c'�G])��� �Yׅ�(�V�Ͼ�)B5��]+�����.({ƥ�� � �au�jk�4����i���(sFA�w߆���lq�`_��+�̢��t6a��sj��h%Cz+�f��X�4B]X�
����)J�>��G�iK��(�ie��H����b�^��L�$ �復j8���*W6�$[����}j9թ������WD��U�X������>L�N٨�kx�Ś�':P�V���|�փ8
3넓���<(c)�����'��Y��j?>�'=gVtæ@D7��s��Q�V�-*��`�L6�Oվ�[2�4�G3�tɱ��*�9
i�_ϨA�5���=��hm���doe�!3�'aJ����Ye �Ӭ�/<�����pٱdB�E�w�}ʃ�idg��2rvZ#�{������Aك���Q�rT�n��'+!{8 !�g����xp�eG�] ��?�	G�\�Q����*}�����a��^��c�|J�y\>�E��&&�Ʉr'�g۱���:����`��?��%�P�v�1�J#L ��L��"+٘�k�� �!n}���du0{o0�-Kn��Bb��B�p6�ܚ��E�4A$�h�_��*���Fs8y�����@�Y���.�uֵ*�evP]�WYS411#g�b�=pH�3�82�j�/�|>������bS�"����s�ͱ���u#�}�w�D��K7S2�+���C��	�XGjy?j��.��P>GO�b�t�)";�Hw�A��Cz"��,	I��I�X{���W&�-ד�H�U��hr��+����X�0/���GD"�&-rU�B�H�^��&˲�e΁I.N���~��{�����9s��Kt<:�m���9tU���m�J� ��D�F�P���p����gt��\�s�i<z��������lAz�5/%*���iz�^����[������~«�{G�[RS	�Ū�a(���[g�D��{�2`�m�0������,��J}�Y�O��*j��}-��aE�U�a	G�P�>�Q�92?����?�U���(��.���#
F�m�s�zp�.���j
I��^=p��LD%?��S��Bk�������D�.ߺ��a�xN����|���H/�-e�Qp�GD59��o�g���&��)!�hH�nӐ����{Ek�̱Eh�F�����&�"��V뀮��Ke������L�I!������u	��|��l�j:^��2�.�I����~Bs$1�Ds�+��#ӥ��Q�N�-���f��;mm�dU�>@�'QON��!��a���uVcUR?9��Eݔ �7W�E��O��(�����[�5��C�sc�9�;��5�h�nʡp-H� Bi*)�m� ����;���{�"���{�r0؎��(���*��gb�8@�.��v񄗮�d��ZR�%���ǀ�^r��B����(��雓������R��ɝ�(�x�	�7�*�&V�,�,\US�SL�R􉛢z.[��L�%s-�����x圁E�'���;���>e�����Iä�Y/%f�.��#�)Յ����2��C5_�
̿S�Rɜ^�%�� w�2��#6��N<F�f�O�<��������J�n'���E`a
؄�tD$?�SOko�4�`�^[aRoQ�D/�uN���xF����tN��"����d��j�('�_B�?S��Ď�����jkT;��B��������}���`&��ЪA�趴���#�B��R ��.�d[���f�]���Z����q�Kq�޵�Cr�I<�Da�F��z���X�g6��J^� ���k�x����7R��h��Ngr\2`NgN������>rk�����
��B��Z2�xF&�t�Qty\D\��QJ����J��[x5P�:]�«�־�|�;��:���dj�4�n4 �S��&u2��D��J�i����~�7�6i2R�`@��^��]�U����Y6��������+G(�.�p�όhl5��zv�c���mQ�.$�p#G^��U��߿[�Ϋ��ŤQ���f�vA)�����'����V��Cu���x>;�}��3�n�+����
���������KHv�	.x�}��T����,�6��*��a�H?�9`��;�D@ț*Vf�,\�ҏ9���A8ȡ�5�V�= �`. �����H��;�-�m)�?)�ޡ�}���iG�En*E����vw$R��@5s�N���P`,A���>���'93Yx%�+�y�B*��C�<�C`�T�d�EJ=P�`�[�:2�J��a�Ķt���3��'[u�:�i&}�}�w��M���(�ն:�!�0��O�G���<����&4����_Ft��q�<��y.H�����c)|`a����(�Dr�����ϼ5����s�
pޡ�
ى���]K�4R�AН֥F�y��j��*WcE&B�	��0�~�mǘ�غ���)s�����1UB�0+Ha5~���s��HҸ��H�¦�c@y����2�%g�X�*��CY%�<N�ո��)V�ӭ��{)(�7�i	��Di#�p�f&����Z�>2w��;����C6b��d!��u�G7�����̀�G�ɚi��Ri|>K�����P/o�{�U�dK���}`����O t9�������dx���3��d����[�]�����r)�)�p1��N;n��޴�O��i�q�*o�����!ÊD[}�훛���zC��!|�kq�%��iĠb�oROA��5�o:���"x,��D��K����?,cO����K���,yŇ|@�+���>���˓�yW�	�Jj�"��9�6���Jg��:}�*�W��,c�x�f����SD�����iΰ��f&GdM���#CD�-��@ \�qESmv��N�t����
� �k�J?�$�5)=���@�����6���ޓ��n���K"ѐe���ak	jP����r�GD{�ځ`�ǜn�A�S��ɟ���j1$Y��(oX���Խ�9>�JK��Q��"�¤~_���1BM�&��mx�[�4�Lv>�-���p>`��Pu#�k��.��Fj�ϥ�]�:�9�U� A�r�Ua����hNYJ�-L�n?�5�E�P��9le����@�,��^�E��[a�C(�� (��ydz�٬�/�$�TG��{�y�4-�a����GK{�T�-�d����Ө"����b !� �F}|S�YfS�PA��Ua�vDU�$ u�iA�lݖ�aS	_%`�WЫ�vk�	r�ԝLB�0;��%�$S6�n5�`G^8\v�+�pvq gL��Uh�]@TO6���Ю �/ms�JIH<#0�Pb�}� +��0~��wϷ�Ґ��<X�os'x"�h���IH���8���p�o>�y�е�G�d%�#/$O�x�!nrȢ"I\1Ou�0�1e�b� �V�|�,�;�Z�F��W��]�����O�~`��	�Fq���ނ~���{<V;�*8�\��J0 ��P�k��e��T?h"!b�İ��r��� �l}����2�T�	����!F�}�o;ߎ����b�u�鷺�W�i�ڎ���HF�b���l%���k�����)rhϘ���=>�	�<wP's����S�_����)�r+e�c����RйR��]�M�u���b9��m*����Η�~kq;bC��_�����P8���N8.�54���P��"����4�pHU3�̂�&t�@�1�٠��,z��,Ry*��U\�
�"	�t��։^8j~��w_N����(f/�6;�@��䳞�������b$�W�)KvF��4�2!�w����蕒4�ݘ��n����N*��
qF9���ń ��tVy���V�d��S�06�(�5�c�����mzH�Ł���*Ϫv���2�,�Ȧ,�69��-@k(D���.9�0��P�0�� �G�[?�Y��u<g�؊�A&���.�W�BM�c0H�O
.3�ZJ\4���2D4Ndlw:U�����l���7{x�7����ݪ,jHA�A��.p��s+��]�B|��om}t�,5�@����������5��eq�����Q����[�{�u��՗��q��7.l�<B�m%��D���M����x�*hH����xz**�c��}G�u8�k�n���gkWp�n�)����_���aᇉ�d��D������w(]��陀��*�M׉l�K�#>(�P�*�ǋ<+$Ӛo��i�n�q�bi��K
H��uە��%O����
b{t�p��6h�Ɨ�ㄩ���J^-h)��cC�$a3j�����H�x��`엚�� !X���w�3�������:�>a����U� ���|!jP�pSx���ś��܊��#�Q�|�I�����?u�>� 4C�BP�]G2M����=ʫ������t��(� Y�@���LYw��l[`)��h ��9^�t���!�xi:}�4�����s�n�6�x���־���Z���^�;��5֡S��B��R�G&�~��(������V�qs23|B�Ů+P�1�R�쥒7�zh�ח���`y~m	�37�4��ӽ���Y����ttNґ	�ēr�B���tW���F�k�/E�+�P���PD�?ʥ�e��辉�`��A�l�Y��t�"F��P�%W	!�ǒ�̶������G�z���
���M���	�f:\����"_�@�r�Ay.������z(5��,�w��ʗT5�
�Z���*��ɀd���[H�����z�2�!�$�a�
"ZR��`������ �qD����;������2��d٧
���������H�����4�5F{�v)E������?N�>]p��R&6�`�-t���w�0}5<6��k����$�lg?�~!M���R��z�!���U��+�������)�;�/��a��OB���L7GUI���?l�פ�r`��L�d\[��6��g���}�$� Co*H�B{�|~F �����3OX^R<b�ݘ���q�	�W�O����C6V�,��O�k�� ��,����B�t~�Y�)�yd�=�x�0��L�l�oN��3�}@���P��<U,��-w���08����x�������]�P�yU�,�t��s�	�2��P���B��A���y'|�`� ���ޑ*���A�?��s���kAݳE?�M�#?�͑H���X��e�{OgSxiݱ4�(�Ej���F(�H�x���'�������3z�il�-����M%�@�:/�7�y*�}"��\�X�i֤I6��ӄ�I(���,��h�LO�"�Z.��M��a޴s�(c�[����p�ۓ9�W��F��rI���#��l�;!�'MF��!��S��,�>;�O=$�f�X��,$�+����m��~ 2����F�[I���O��Y	�s���0�23�`X��E\A?�{s0�l����6��JU#���b\��S|q�������*�����X���K��2�P�Cʸ �;����A؆���Vx~��&ԟ{>��:�t��ۍ��O��%���]�g�v�����"�_r����7��%��pp��<
�����n����j���`���mD��7�*�#���ʝ�z*���I�Crl,�!q�j��P�l�)��=}��KN,<"E�A�{	Q?��k�T��5��'�0�6�#��Z�P��`Wq�H�����y���)sv͍�
����bw�V�Jn���s��pꃌj�gV@X���N��_]3��������і)�iTD[Tz�*�2cs%Ȩ6B���A�, ��k�zP�*�6@K��:5��O��u�F�y:J�ُ�B_�j��P�O�]�/��o�!MG��m��W�S,���O&��eԉ�Y����6�]��R�?!P4�Ԗ�NS��Z|񡉽��5D�X-�ߚC~F}
 3`2о]��V�8	"$�ĶJk�w8�<cLH�:%�Kj�M]�`�&;�R��~�![]�0DZf��ӂk�n	�L�$	tWͲ�2��fK�i�'ACb%_.���]E�NrzCW �w����oߝ?9n{J_��N��`�_��7/��c��㜋�J��kh�Z��G������Ļ��ŗ8��u5���%*���-����r'�����
��`O9�u�iXK<NO�_^������E����!�I0��}�C��6��>��p;\4?�c���c�P��f��/�Z5M��=�F�'dh���I+$��니|Z,ih!�Z�����mՏ��ܝ���yrY�P8m�~�x����b������FaMk�.����2U�M��Ĝ>�H�vr��o�|���kd�q��9���v<yѵ,~_�`�NXA5P�L�+�N� |������R�GLH�Ws3�	�Db���*���a�4n��@��Y��}�S8֍�i���:�]�Ž�AN?gToV2��͚�:d7���h�9Zg�8�sm0�\ʅ�J��yL�������J�t}i����n�R��@S��V�Д����h[`~
��)��W���	h+��8�rKVC�`9��|ء���a�ހ����r��5�@OPW���������1����U-��))QN�Y�x�4&�Sx�&�Ium�+��^�ӊy�d°��Xr��cK�~����8(_K�+��TJ���;���-;�5��h�&�y�n�{��� ���@�b�ז�`�1sH���&�Y��6�E���Z���� U����WdqSG���7>2�px�����,��p��0E�;k�,M���p����A����-<�4�J���=�=Y
�I� �!��zF1G��O�&��ͥ��ϱ|a�2�ԁ6[���\�� (p�w� =N-z�,��%U�hE��wg��qX6(�H��p���ˠ�w��&DBӰI�(��f]��G�S9I���b���V}�������ߪ�;^���->v�S>`6&�+�%���c��Z��a�8�x�@�H`�r(�~EF[K�;�F��DYG�`�	�2|�nmҺ8�PhC�D ]O��\�V|y���jILRN'<'�g�A��{\({��mX��%�\��/�>�a��/�D{�=E�Ś�TC��<���Bh��-��7XwV�kG}49��;9����,��?��\�h��x2��FD:�ܻ~�~,���T�M��6½���`����{@�~�(j��K�$��aRt�W�_�+�ql���Ș K���(V
��JhU��b�i4(\�ߗR�2�m,D�L�\�� ������8��cЉ�?^��D\:6��u%YO���go��Z�T�)ulAU��kp�0����)E��5�D ��6=q��]vx�lk&��d��l�jʹn�	��S�V�i�E��f1Z굪 ���S�w��E錏��%J� ���Z:�9�nl��=P�Zd�q�h�[�hgn�ERA�Y�)��GrC�ћ��s��g6ÃB�[@-x~{��+�`�0%��T����hހʓJ?vv:Į�«Cj�!����[���cCX�F�P} ���
ٷ���r�A��!�u�O�<�2Y�jJ<�x���v�b�Ik	L~�uU�D�k?���1�@o.zYڰ��v{dL#)%~���M�U�e8�^�&��K"��b�JK�	.)��'~�m�Β\���@����Eσ� sZK�dЅ�����<�~���8?2�~�_>e9rsI�i# 4��|��C7��e�b\[u|of<#��&ǜF���J�UH����6�ڹ�6�(�=�މ/I�����9�{��9M���B�8��":�|�d�)��I	ו��(/U���y��'�a��Ό<���A��J������l8!)�"g�e���D"0�ƭZ���;��B�2,vX�+n)���	�FĴW�<�%!�~8s)'M�p�>�b��-?�T�'b���!'���a�Y�8��᷈�m5��d;�����A,���p�Z}[\4%����H�D��.:�mJ�7=%(�$�iov�����iKN�Ǐ�r�?]��"S��~T�����&�����ѵ�˕%D�b��%5��-(ʒ�(g��ge�:�hm��@�!:3�!z�h�*0�t��5��U�����a_s��Bp�������DQ��rfU�"� �*/{B�ҞQ�FZ���zD����O���HnX�]��_z��O*P���:�D6#���%� ⢃�cx�X���������NWa��ڂ7(a�'DhƍXE/T��^`�K��
r7��n�z�x
�[��f#{*@�Wa�Fd��c�'�r�{��f�Hf�@�Wc@��Ԗ,C�	�	�F@�u��8��r)�k`���ATg���@��F�83m~�S�:*cX�|�_�_@�Z�(��K�㛩��pm����^�`��}��܂�QJ�K'@�4_�W��U1�a��[vD��X�D*�����lռL3�.U`��,vy}��w�s�������82�n!A��-�@kQ���z׷�G^���Ń�z3z"�,d#��z�P����_���`*��m�^�>�v$��2U@Y�'�� ,����F���� 4�������q�u6N�����l��?1����Mp(��v�bݎ�/F�a0żÐ!����g��X���;�'��!��|�s�a	J�4{_mH��䗒�f��C㮿i��ǽ�9"݄��vc�P�㺃���*��t��b��6T˖g��ݾx��v�gYt^���BK�Є�v>2��P�������P؝ ���W��ņ�_��XM4�t�*�7g���[�svH޵jS�@�!w^��,�r�plD�/��<}M5�$�{�@$�[P��룧���_�r��M��R��D�8��K�o��_��G}Di�-����>;忈T����Q}�`F�W)كI��^�	b�s)�\N��-@��	�>�:��9��4��Ә^'��	14���8�ek�@8���뷞	XM|Kc���3�i�f9�R��7���7l6���Qk_�\���3���#��$㷟x�T���
ߎ�P�d�c��`�Ieq�������2��h�3��Jh���9+�i�)��h֜�t�
�r�1>�!ʎ��CB�{��G�6A( /V��G���ҙ�����#[s?8x��/�"iX��k?"��sb���~�����H�J!�փ�-4�*�  p�!>U�Jlhb��4����� �I<�H_�Ѷh$5��
��Θz��늈���J���<Rפ��A���"��Q���9��n���mc�;���iG�90P�X�îf<�o�52#�I�f�y��M�wH����J��J���|/5h����X?|RC��c�@����c�׭n~���vv��?����X���R{G�d�c�1���_K�s^����67�?�˷��Ò��'�	Vݝ�sy��a��D��N-�D�n2�T�ΰJ3�\p�*��"�1�/�هs9���A=d��g�4�_5;�O;t�;�^<�gj��(�np�d��(���'�8lC�E}�hV^���:�>Q�fK�ph6e*��S��;;2�*�[���|��s�h:.]T��I�L���e1���D{�y�Va�*���a��NZ������zìz�g��!�-P��M��%3�j�2a-���ܝ��er?��V��&�v��6{��@�=��xٴ??O��:V�T�[�YE�p�LUw�qy�&�������}�����>���#B��ܨnkdH-&}Yo�N���h�S�iR$�9�B������m9�fF��i��kMv��5���'�%*3Be�H4e�끋|eJ)��SO�_i	��d�x���?�\�L�3�-d��Z��#�5Bg�x Da#;c�v"r�pD��{e���XF|�`3��Sv̗��_�F5W]c5�i�p�W�5 /�K%o�	4!o=;���߶�B�@�%ňK���Z��r+֯u*( �=	$�#G��Q�H�h`m�uLJX3z%��Fo����b�I��u�J��]�l�-U�D�]���������QXPs���y�xm�Ѻ&��ۘ�K�Rh!�� v�\��<9_u� c�6�x1�屈�CI�:���t���g�q �:�R ��k���Ϣ�Kj�4�ŋ��P�E�l��H���V6���c���r!�.����d��Ѭ�o.j{6��R"d2���g��<�yٚw�^J�ն�Nt�z;~�6g/��[S����/A��Ι���r�T�%^�E�S�C�IW���جg���|y
Ⱥ�NT����Q~�����8c������a��]�~�~Y�z�{�`�9�NH�O����3GHˉ�D꽴�c�<�wsnw�)Й���؊oA1�����6���S������ "=��Y,GCe�,itƿr����8WEǱ ���(�o��ZјS���@l������`�Qa	֬aJC�L��e�f&Gި�	ӕ�?�h��	��D�0U�]�����~��_��e4_~�����!�5b�5=�,���2=���e�-=��bN�e�R �u��VkH��׿p'�+�]��b/�ƨb$���v�-�RRy0%�z�>���5m��q2��`�%�D ��SQX�:��ӧ#�~N<4YN�|�A��LI�M�w���R=h�smp��E��B�m�
I��r��K�:42��+�¿~S�r����
p)cb@�;�ٹ�Į	���v��5�(�V|��f�^ i,;�Ʉ�����ǢA&��wZ� ~�]�����C3۝qك!2 ��Wf%��N�z��`���Ui���u٤˻�M^�(`���P�]�﷾��y�?���HN�<��$�8k�&�����~�����	ˮ�s�
�o��]�E?\p� �X�<�OI];�BG~A�-���r�`��:�I�ͷ}k�|pp�\�` I7RqJ��;��\��OL3`����冰k�@]J����"&.�U� �M���*�t���ڛZ*W����D?������l�G�i�*'�q�@򶫻S�Bd�C���[m�����ef|�H����ѥ�-i�2�';�C�d3f2�������|����Ĭ�n�F�QK�1 <��.p�B�y�dR���N�װ-M�'Zc"�A5ڄ�ҷf����U�-���w�}�����U�����^a�a>{	�pJ;�/h{�=�{m-�غ�T��%�C8b��Y6)�8�jT%�?��T�"�p.�9b�v�'��zS���a�L���6�b�B h�F���
�.7['���5����l�W��'��_myAɜ�.T*E��0�i|\���3mlڱ���x�HU=���Q��;L����8�*eq��˄ڂ�<<7�>���Ϣur�Vw�~�U9i��]�i�M#h�}�JٌP����~�N�)U�`�-���Z�QV�+C'�/��[�&p�<M�%F?pV'��X���\謯�E��"6f �o�2��6��5ɟ`�j�Y�R]<!��b�&c\`YHCG�;����� I�z�T����|���[��Q �w�� L�£��z_p�,��J	����y�Lf�{���ϫ�h�Z�?W^�׌2ټrLPȷ(�yHQ{<�^U0�ca��+!@��9Kl8i����v�
�+n8h����;f$&����5(���G���k�Zes� Qx��gZW�ȟC��1���