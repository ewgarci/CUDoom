  --Example instantiation for system 'new_doom'
  new_doom_inst : new_doom
    port map(
      SRAM_ADDR_from_the_skygen_0 => SRAM_ADDR_from_the_skygen_0,
      SRAM_CE_N_from_the_skygen_0 => SRAM_CE_N_from_the_skygen_0,
      SRAM_DQ_to_and_from_the_skygen_0 => SRAM_DQ_to_and_from_the_skygen_0,
      SRAM_LB_N_from_the_skygen_0 => SRAM_LB_N_from_the_skygen_0,
      SRAM_OE_N_from_the_skygen_0 => SRAM_OE_N_from_the_skygen_0,
      SRAM_UB_N_from_the_skygen_0 => SRAM_UB_N_from_the_skygen_0,
      SRAM_WE_N_from_the_skygen_0 => SRAM_WE_N_from_the_skygen_0,
      Sky_pixel_from_the_skygen_0 => Sky_pixel_from_the_skygen_0,
      Sram_mux_out_from_the_skygen_0 => Sram_mux_out_from_the_skygen_0,
      ctrl_from_the_niosInterface_1_0 => ctrl_from_the_niosInterface_1_0,
      nios_data_from_the_niosInterface_1_0 => nios_data_from_the_niosInterface_1_0,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      Cur_Row_in_to_the_skygen_0 => Cur_Row_in_to_the_skygen_0,
      FB_angle_in_to_the_skygen_0 => FB_angle_in_to_the_skygen_0,
      PS2_Clk_to_the_de2_ps2_0 => PS2_Clk_to_the_de2_ps2_0,
      PS2_Data_to_the_de2_ps2_0 => PS2_Data_to_the_de2_ps2_0,
      clk_0 => clk_0,
      hardware_data_to_the_niosInterface_1_0 => hardware_data_to_the_niosInterface_1_0,
      reset_n => reset_n
    );


