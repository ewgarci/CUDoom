-- megafunction wizard: %FIR Filter 2D v12.1%
-- GENERATION: DEFERRED
-- synthesis translate_off

ENTITY anti_alias IS 
	PORT (
		clock	:  IN STD_LOGIC;
		reset	:  IN STD_LOGIC;
		din_ready	:  OUT STD_LOGIC;
		din_valid	:  IN STD_LOGIC;
		din_data	:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		din_startofpacket	:  IN STD_LOGIC;
		din_endofpacket	:  IN STD_LOGIC;
		dout_ready	:  IN STD_LOGIC;
		dout_valid	:  OUT STD_LOGIC;
		dout_data	:  OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		dout_startofpacket	:  OUT STD_LOGIC;
		dout_endofpacket	:  OUT STD_LOGIC;
	);
END anti_alias;
-- synthesis translate_on
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2013 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="alt_vip_fir" version="12.1" >
-- Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
-- Retrieval info: 	<generic name="PARAMETERISATION" value="&lt;firParams&gt;&lt;FIR_NAME&gt;finite_impulse_response&lt;/FIR_NAME&gt;&lt;FIR_WIDTH&gt;640&lt;/FIR_WIDTH&gt;&lt;FIR_CHANNELS_IN_SEQ&gt;3&lt;/FIR_CHANNELS_IN_SEQ&gt;&lt;FIR_INPUT_OUTPUT_DATATYPES&gt;&lt;IODT_INPUT_BPS&gt;8&lt;/IODT_INPUT_BPS&gt;&lt;IODT_OUTPUT_BPS&gt;8&lt;/IODT_OUTPUT_BPS&gt;&lt;IODT_INPUT_DATA_TYPE&gt;DATA_TYPE_UNSIGNED&lt;/IODT_INPUT_DATA_TYPE&gt;&lt;IODT_OUTPUT_DATA_TYPE&gt;DATA_TYPE_UNSIGNED&lt;/IODT_OUTPUT_DATA_TYPE&gt;&lt;IODT_USE_INPUT_GUARD_BANDS&gt;false&lt;/IODT_USE_INPUT_GUARD_BANDS&gt;&lt;IODT_INPUT_GUARD_MIN&gt;0&lt;/IODT_INPUT_GUARD_MIN&gt;&lt;IODT_INPUT_GUARD_MAX&gt;255&lt;/IODT_INPUT_GUARD_MAX&gt;&lt;IODT_USE_OUTPUT_GUARD_BANDS&gt;false&lt;/IODT_USE_OUTPUT_GUARD_BANDS&gt;&lt;IODT_OUTPUT_GUARD_MIN&gt;0&lt;/IODT_OUTPUT_GUARD_MIN&gt;&lt;IODT_OUTPUT_GUARD_MAX&gt;255&lt;/IODT_OUTPUT_GUARD_MAX&gt;&lt;/FIR_INPUT_OUTPUT_DATATYPES&gt;&lt;FIR_FILTER_SIZE&gt;3&lt;/FIR_FILTER_SIZE&gt;&lt;FIR_SYMMETRIC_MODE&gt;true&lt;/FIR_SYMMETRIC_MODE&gt;&lt;FIR_COEFFS_MODEL&gt;SIMPLE_SMOOTHING&lt;/FIR_COEFFS_MODEL&gt;&lt;FIR_COEFFS&gt;&lt;kRow&gt; &lt;k&gt;-0.25&lt;/k&gt;&lt;k&gt;-0.25&lt;/k&gt;&lt;k&gt;-0.25&lt;/k&gt; &lt;/kRow&gt;&lt;kRow&gt; &lt;k&gt;-0.25&lt;/k&gt;&lt;k&gt;2.0&lt;/k&gt;&lt;k&gt;-0.25&lt;/k&gt; &lt;/kRow&gt;&lt;kRow&gt; &lt;k&gt;-0.25&lt;/k&gt;&lt;k&gt;-0.25&lt;/k&gt;&lt;k&gt;-0.25&lt;/k&gt; &lt;/kRow&gt;&lt;/FIR_COEFFS&gt;&lt;FIR_COEFFS_PRECISION&gt;&lt;CPC_INTEGER_BITS&gt;0&lt;/CPC_INTEGER_BITS&gt;&lt;CPC_FRACTION_BITS&gt;6&lt;/CPC_FRACTION_BITS&gt;&lt;CPC_COEFFS_SIGNED&gt;false&lt;/CPC_COEFFS_SIGNED&gt;&lt;/FIR_COEFFS_PRECISION&gt;&lt;FIR_OUTPUT_CONVERSION&gt;&lt;ODTC_SCALE&gt;0&lt;/ODTC_SCALE&gt;&lt;ODTC_FIXEDPOINT_TO_INTEGER&gt;FRACTION_BITS_ROUND_HALF_UP&lt;/ODTC_FIXEDPOINT_TO_INTEGER&gt;&lt;ODTC_CONVERT_SIGNED_TO_UNSIGNED&gt;CONVERT_TO_UNSIGNED_SATURATE&lt;/ODTC_CONVERT_SIGNED_TO_UNSIGNED&gt;&lt;/FIR_OUTPUT_CONVERSION&gt;&lt;FIR_CONTROL_PORT&gt;false&lt;/FIR_CONTROL_PORT&gt;&lt;/firParams&gt;" />
-- Retrieval info: </instance>
