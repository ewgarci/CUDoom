// de2_ps2_0.v

// Generated using ACDS version 12.1 177 at 2013.05.02.00:39:21

`timescale 1 ps / 1 ps
module de2_ps2_0 (
		input  wire       clk,        //          clock.clk
		input  wire       reset,      //          reset.reset
		input  wire [0:0] address,    // avalon_slave_0.address
		input  wire       read,       //               .read
		input  wire       chipselect, //               .chipselect
		output wire [7:0] readdata,   //               .readdata
		input  wire       PS2_Clk,    //    conduit_end.export
		input  wire       PS2_Data    //               .export
	);

	de2_ps2 de2_ps2_0_inst (
		.clk        (clk),        //          clock.clk
		.reset      (reset),      //          reset.reset
		.address    (address),    // avalon_slave_0.address
		.read       (read),       //               .read
		.chipselect (chipselect), //               .chipselect
		.readdata   (readdata),   //               .readdata
		.PS2_Clk    (PS2_Clk),    //    conduit_end.export
		.PS2_Data   (PS2_Data)    //               .export
	);

endmodule
