// skygen_0.v

// Generated using ACDS version 12.1 177 at 2013.05.02.00:39:16

`timescale 1 ps / 1 ps
module skygen_0 (
		input  wire        clk,          //          clock.clk
		input  wire        reset_n,      //               .reset_n
		input  wire        read,         // avalon_slave_0.read
		input  wire        write,        //               .write
		input  wire        chipselect,   //               .chipselect
		input  wire [17:0] address,      //               .address
		output wire [15:0] readdata,     //               .readdata
		input  wire [15:0] writedata,    //               .writedata
		input  wire [1:0]  byteenable,   //               .byteenable
		inout  wire [15:0] SRAM_DQ,      //    conduit_end.export
		output wire [17:0] SRAM_ADDR,    //               .export
		output wire        SRAM_UB_N,    //               .export
		output wire        SRAM_LB_N,    //               .export
		output wire        SRAM_WE_N,    //               .export
		output wire        SRAM_CE_N,    //               .export
		output wire        SRAM_OE_N,    //               .export
		input  wire [9:0]  Cur_Row_in,   //               .export
		input  wire [9:0]  FB_angle_in,  //               .export
		output wire [7:0]  Sky_pixel,    //               .export
		output wire        Sram_mux_out  //               .export
	);

	skygen skygen_0_inst (
		.clk          (clk),          //          clock.clk
		.reset_n      (reset_n),      //               .reset_n
		.read         (read),         // avalon_slave_0.read
		.write        (write),        //               .write
		.chipselect   (chipselect),   //               .chipselect
		.address      (address),      //               .address
		.readdata     (readdata),     //               .readdata
		.writedata    (writedata),    //               .writedata
		.byteenable   (byteenable),   //               .byteenable
		.SRAM_DQ      (SRAM_DQ),      //    conduit_end.export
		.SRAM_ADDR    (SRAM_ADDR),    //               .export
		.SRAM_UB_N    (SRAM_UB_N),    //               .export
		.SRAM_LB_N    (SRAM_LB_N),    //               .export
		.SRAM_WE_N    (SRAM_WE_N),    //               .export
		.SRAM_CE_N    (SRAM_CE_N),    //               .export
		.SRAM_OE_N    (SRAM_OE_N),    //               .export
		.Cur_Row_in   (Cur_Row_in),   //               .export
		.FB_angle_in  (FB_angle_in),  //               .export
		.Sky_pixel    (Sky_pixel),    //               .export
		.Sram_mux_out (Sram_mux_out)  //               .export
	);

endmodule
